PK   sRWZ'.Ǐ�  {�     cirkitFile.json�]Ys�F�+)�@���6��*?d�J�������.EjA�N�����q-u[�l��f���i4�/A�~*��|Ӕ�Oe��7����Ep�6����l<��e�Y~l������<�a�yxܬ�u��e')�ì�I��̄	�EXX&�TLf�-Yp��n�bv�c8v�cW8v��ǘ����8f�m�jm�<S"3*�m���gy�cO&.<��J�R�yg�r�B�<K�sS��!��Nh�VT�,d�t�B��lgL�0�)gڍ�L�4s�Zm���Q�5J7r�r9a{e
Y�B;�8��<fa�ıCU�L�R��Mrs��G�R�ܦ|j���^���"�2,	l\B�^ #�@BW �+:(G+��(Գ`T3(�L���"CMr�I�n���&�i r�H�n�HG/���Ho#�I~P�1X��c��}z�@����O�!�J��WEX��5Yh3�
�g:&.X5�gA��<<H�i�F;�	�i_	+�H�_��a�H�wI5���=�[��(���,���$�.B��:xB�H��i��/��&�C��]@��(L-0!4Om`��-����Pm1��w��-�X�C�Fi����t�oV�Y:�g����ZA'�"H�H)�D��R,/X�!�[b)������!�z)���mC\9;�^!�s@/�Ja����w�ʹ�U�C`�i��@��`�w ��I�ci��D>�ł���U�C�b�Ј�A��A��A�$J%h�'i�'i��������r���-��Y�Ak�Rf�Z�%�2�_h�����^	l�Aݬ�Wc)�Рw>��h)Ĩ�\t������s�Z�����5�o'h���9�PCk��O>����y������G �ϝ��ն�@�nR�\Z;�r.�m۴-�%�u�k�t�,��)�D�"��I�)1���D��Axi��i��i��i �i�i �i0�i@�iP,hP,�|0��������%�%�%Q*A?I?I?I?I���,��%1��Y��Kbx)��.����\�K�E/�$��2�:�%114�Oc�%114 �Oc�%��b�%1�������Rf\�*\�K��]pI/�Ɩٕ���Rf�\;J��p/o�=b˺�=��j|��r�|\�yY,��r�e�|��\b�y��|y �'4c�c�=�|3u^è��F5�5KN��F\TE�[��x(��mT{.&�|��@b~V S?~+͓�ɿ�5�B�����}w�M����x�.��g�E�;�|ʀ��Wx��� ��`#>�l�j����i �	�l���|;���u��
)Bg ��^��W��30�^#c�^���Zf��5l����2 t9\��z}jX:��T�&:�ʹ�l/��ń�H~��WH~_$g��o��91�?^΄K�,]J��e��y�����ӓcۙP�IB%vXxw7�P���XH�L��u�uyX�+�N�S�u�L�fטԃ�,+�8#8�&%Th��Tbq*��f3���+�ݫ]�ф p���
���E�+n(���䘘����~�suXt]qs�V"� ,>�����!� N��C���Dԓ7q�w�B-���J���&V�Y�3g"����M�I��F0�n:�I�p���#2�mH=�0_���p'���-I=q����.�3_]����E.H��x�O���6�=�=d�K�nȻoh��SrO�=mw/���������{�9���l�!<���s�!<Gw@x�9�琝9�Xzb鉥'�^��~��I���8�q���G�̎��Km^ >=&��=���Y�Ln�+P?M��.�E��a�&���a������޷a�D=^ �7���L ;�)"�i!Ȧ�a��{���n��➜�k������z��	�g�qmYÔ���}�s�j}'�*�ʕV=}������k��Ð�Ð�Ð�Ð�ÐŇ�x8����Pw�َc#C�0d}���Vˬ)�"ۤ��o�6�U�m��~z�X��6u�}�>z�l˦��.�|x\����:�۶���=��������S���w?�����ݺvJ�j{������NnpS��m��e�[���Uy��)�����n�fW��zH׻*��]S6�xJ�Ē���6-�%�W36ۺ���Ai��l��Z�Z*���/qs��|�x��(�Ը���4㠯����UR�R�������vz�"p�~��� PB�6M�{;�ݣ�]7��<��%�H/�dw��k�DLj'��~(����6fz!��!�=^�r��(�2�|�@�ȉT�N��8�VY�L���Ǣ��P���N���F�`Rz�U���<�������<��|��mF��BX�Ds%�a�{���q.&��Rhwa,�n�����7`�^�H�bϡ���e�ȕ���|:p�-����vWԛ��H:/1��/�-�E�]�_x����O!m�l�,*w�����(Y��IÔg�t3_�n��Ct�@Z$�J�y�LD2V�E��w*:�G�8*I�%�����n�K���qT�J�%�l���E�����oEZ5����ݺ�yw!�ޔ�XDF��-��k�V�8�O��R˪��NY��
�M�����*�,tV Ϫ�/=�V�;���a�$w"�N�sC�y���Q'o�d�*�|�Hì�R��05i��)��R��Ԡ)U' S�Yc��sęeǗ\?�� }� �__a�@��1?����vzi���'(��:�o.��Ew���������,U��C�V�
�C�biX�<)La%OaY�P	�����OGhb��V�Ǖ�l�ʉr���}c�:Q�#�<�{�F��t�6._(#���9��xl@d&���%0i$����IS0i&-�IK`�6XS�/��蒎RVt�j���T���,��p5G��9J5X�Q��R�RVr�j��cT	��J8H��h�P�8�@�8�\��I�H'HSd��Y6�����`�K�ݺ���v��� 4��:vVe�SO�.҇?�E{�>6���u��}Y����;�H0�q���vK�����T1yߔm��ou����ۄ�L��6�~-�6��=���m��uyuڴ�����z��NX�.����`�D5��_)Ms��Ag��^����������6�����~�����|��v�6;�-/�nO���E����;F�ET]���\�����z|u�C�x��m-8~�c @�0� �����p^���Ǡѕ�ЀQ)����/���7��3�{h�s�آ�O��U��S�_�[�o�g���~c�u}2ia�c����0tA�S�Ð�p\�f��ѧ����Q]ֱ�T��uh�?@	N�oHbhp�|C����)h����N�/�ŝ
 4��?T�����E^�R��,��F�J���/�L�V� ������l��R�1�3'����9�=hE�I����!ˋ�0�J�B�|\é����
����H�FX��Ϩ�<�82���:sYG�Z�����N���T��Є�0��д�0/ʃ4}�	�pj���].����?D����B}x��U����8�g����9��e���Di���&Vp�uH�5�y�g8�g�F�^����h�ҧ�A�W�R;����#�(�ae�����^�.�O���ؙ˼F6U��wD����꧴-�:]m���m���Y���w���û�|��K��zl6�)���r�7�㡹&��'PK   sRWZx^��6� _� /   images/00531496-7d3e-47f9-840c-8f79a4e99c6a.png�e[U�7�	%AJ$EZZ锖��t�tw��t*H� ��i��nx��?�|����.V�9���k,��*Haac�`0,�7��0�vo�>�I��	9�����{}#=_-�?|�,��bg��f������bak�dlh�����,uG�{�QuOۚqsW����~�{��SG��A#��)��C"�9��-���LY�YY%�o4��k05^�4աs��2i�=K61x��������S��<=�����*�����f��fz��%����#�m�A�����{���=���(@��#L��{|��E�]��4[���0����9������C[J�P�>����O�i�<~��@��X�	%%�[�{777����		�S�b���9_f:��/lMTt����S���Ow� �BQ$ܒoޠ�������EECC�̯�q&���y?j)���^�Sk�����x�?���i����N��#�5[�g�`�s��Z��BC��P�<W�����fFF>L�s������|����0߂D�s7M����b��9f�*�
Ӿ��[��X�����VR��e�e�]�Y�$9Z��3DVֳvs�n3.O������Z�9�d��ikC9o��č���nO~�MdU�e�[=8%�+����)8i����2����	aĽ���7o޴4�\�UUU��?{�3d.��}��ܠ!!a��L}�l"KhDDaUP� �S�{����hU�3�׻~�d�P��\����L�/�ʕ}2�:e3J�Q�����x\�����z�� �E��}ϙb���X�l>pm��Ivv6�?�������l�Sn��8*)?�]�%���H'Fl������#���B(@��f(=8iׄ^+�O{�6�_�w9��VB��]54���g��.��d``Шwe沙���~q)t�F��`��(���g���ѽz5R����?����,{�KX�[O�u��!^n�	�3�Z��C"6���951����>#33VAA��~o�+��y�݉^��j��
TЎ7FŮ/��~X�}���b���w��?>�Y8�^Q�?��o8���x�la��Ak�MB����/b!�n��ܕ�,+���x<�����).M�:����8m�ɣ� �p��S�{���\���顡�!:6v�v�\4��ƴ�7l�r��x�W�F�� ����PfR���(�;�K���͐���M_?SSڏ?p�ƥ�E��<�l�|~�җ�9������%ayy9���V0�
ߖ.
?�P��׻%���K%��+���|p�_ϧ722��ʸ'�s19R1�eee�5�:��pFq))*pM�O=�:�5��/�n����*1555�8v�;�1 O��2jJ,����\Ɨ'��|�����S8��Yt��3�vD�]�K6�>*ߍL���a�]I...�mUd�\��71mMV>�w�j9ٞ���YM�ZZ��kkk�:����t�x���q�Wx�jE-xa�O*�<�i������ٶ���͑��l쪚h[�K�o�����H���/�F�a�`	���1��bE�V��m�!a��B�U��<2G�J�ɮ��~�������p ����^�"�]6�f��\"H(�Z�hj�Zfu_�M��m<U;K��ʆ�����UGG����mN�Ѵ{�"�Q��l��o����?��c��c�c����֔A5�Q�W�B����K���ݩY�ƼM[__�hpgo:[|�Q�2����h�=-�������c��1����j��2�ς�R�����ܖ��]�����D
�ri}�6>��R+E�?
�ӧ�_v�C�{�'��ӡ�"��U�X��b=o���"�=��=
Z�iq�~s�o�%����z�-�X�J-f�G�<����U6ڷ���`�p�s��a��{N� @9�;k� ���:]�9�wu-%�������9c�6x8ɥraV�0y{�Y�Q�HSe7��LyC���M��<�S������ Dn<(���D^Cm��z�SQ���dCX8�����������YaQ
tt?UW*�kt�ZY^^H�kj�f�؎��w�/�A��~࣬<|#�u��������8!7�|E�-�$LH}��n�������vԙ6���R��B`qK�F �����̪��m�;�i0�^=��YV%��)�����McG�4J�%pg���Tc�Ï�f�D7��p�����2�­�A �rOu�V�xz�脱6����=�5�z+�}[v3�h[[��c�������u��=������;�gBB� Ylh�6|@�����!H�������j�_g�D�͊�݀�I^NN�8\�P&��F4"<<�Rf�y�9S��n���!�@�4��@f�fis4�t1�'4b�)l�䗹�T=���{��Wh�]8a���ư�Ĵ4�/}����G���=j��_:���kW3�@��O�:��*fDF<aU������rJ�c9�1F~�ލu�?=bO�D?<���Z��j�Gǿ�ᰳ��m�S�+�h���?k�-F�B��nG� ���f<�-A0�	�{{6=�mΣ��߮��� ��f|8l�;���=ӊ�qD8�\�'C6�?SH�3$R�]5���	�^;@�r ���9�"nN��ZH��v� �$qۑs���x��O����KD�2sq�(���({�o-/�����ç=V���F}�J�p4,;���sW���n�ᣟmm�֧���PP�b(X}������M��Tʠ�r�*��OH?\Lو���_\nU��N��+�0���G2;V
0
��L� I���39�2��=�� B��U8z�a4�4Z^���6�6o�mK�������^g�a�z���W�c���;@��TZXK��D��H��A�� �u؝ ��K����2�����6=���x��)�滕�>w$���Lʪ/ �mxsu��č�ad�Ê	�l=��A����2]m�W���~��[I��؈eN[G'R���p{�NJs��P�vF���e���v�䒶]cn%�4!E���7M��А��x'�������n�{@��޷�#y��N�s~�o��� ��;���|?��pGJn��r>)^�g��u��s��>��S����(�S��>��n�]��^�����]��TЁ�d�c�H�2�|t�z��;�p����.@�u�[?|Vz��_O��ݕ����K�ց߿ۃ0����E]��g~w�Q�_�O�e��'H�	(��c�&�dQ�]���fj��ŋ�\�G�F�1��� Q�})�޻��S� N��w3����S�)���h�0H�LN����`f�jDo�***� "��t�GP���lzY؏�щ�=�rI0??��SÃ=g;��G��̠V����; ���	�nu�P�{^H��?���0b�L@����֋4���"7�w{�2���� zz���g�᮴�D����ϧO�+���0K$/�(El�F��
<z���y}V�f��Ͽ�~u~8�U��T�aL�n�b@h�A��u�r�c��`�˔���{`	Ys�c�ddd���	��~��T�'�I!��q,f� vh·G�	� ���*3��M�
 x��x�w��A/+Yan����֖:������{��ƳDP�4�` yRv㔍v�k5*-�� M�HȻ�w�eL���8�
��>!;<22A�/�V� �ǿ�r�|�������)Ґw�)Ԯf�̬��w����d$�iP<M�!W����'��XP��`d���suF>]����=�K����>#��#p�L8Hu�|����α�´?-��i��v�C�WH��������|����}��s�]M���!��sxO�� 8�Y�RP�g{mغ����(
��x�J�e�iW�;����A�((�Sa�0z&�v��F5Sd!ß�G�㊥lҁQY1���@
�4�Vj�{�X�-kգ�m�������Yj	�3�ZVT1P�ͷM�K� �#+;���q�J�$�7�Cl�r)��|�2<���kGJ.����`�0���+$��2����0�����B�R�?:K�������j�x���jP��7�H�{��V]����w�|`\L�$#��ƴh�3� �mPxyD�w���ᐜF�����rjN�zU�W����n�NR�
�MB���❜!Qoo����p�{��pJ�y�)��b�> ���x98���b���w��B9C9���k��/|1����0dX����;�c��׼<�&3���z�\"�T��&j�X��ϊN1� ����{]��(XOUk$�|B;���؜Q�S,�aJ�w+1����]m�ߊ��cƕ쇡
��[�d���c��'��ODC�$s�o���"<;�e�J�l�"#I)su,���I���X&p^�&���S`�Ȫ���
���d�-���4���.�R4����������jՖ�/no.S��DE�f�v)yx4��z�p�� �£��L����;'��,oT�Hqmf�^z������nW���[��?zJ����Ǘ�FC��z-G����WPT��Wʱߙ��J�?���?6,�P ~l��ژ���I�*�4B~e��ރ�%\�Tqp�}	K\R�R���'EHHu�o�f��0F����r夥�b��Z�```$�|�����'�ݞ�w�L�TO�w���ӊ�����½4��rOS�_�3���44�J�J4ak���}`uRM/���a��2
d��bx�5��wSŘ�M}���Ic^��P���MY��/�e*}�/ڂp6m\ >b�cJJBb���f!��^d� �De�^0����;�P�E#���-&���p�%r���K���2�[߾��SR#c��Cf6䄄��z^��K]��~�w׿T�����G�W���.on��ύ��v������Ж%���;��`�|m��b�2F���=C���v&��H�*�� gQ	v�������}Ӂ���5��_��J��Y[[֑$��T߽�p��L����t �777װ4�!�t.�h2��?j��-F�}�����K.���bƳ3�H��	�s�$c����haq�Kr�J1L����K��qx6RR��!������e�2~d�J�������xG�^7
���T��BlU@���yUX���Hм��@~&��9�d���cc�&�u/hº��#PQ���^�h��}ߨ�
�'���c�>:� rb�pv�Ns�ˍ�R ��<j>q?�gy��A��35���/�����S';3$�3n�
qН�,Ă���ƫ4���)Hxz��z�K���3p��-���[u0�+���EU��w�yuꔥ��y��YY��. �ן��t*�AH����&T� |{�tu4��b����"M��A��R��� ��N�D�T�hh �I��J�2o���>��Hg�c'�{����g�)����k<C�^5��v��ym^�5��h}$.5ժ���'�������i�/	j.�����ׯ���bHF�� �r�Q>�����
�t
i-��MV�(]X�n0�ls��`P/Nz�2�m�H�f;��Fl`�;x�z�3���U7�~�^'[E��\�#4lu�@�h˜s��`5 l�9�[�������ۨ =i&-Um;�����n�D.��W�954�T��r혝��(l�K�2�6 Se,���J�<| �b����t�Y���KG~w!8?o\�;��n.�,ڂ^o��e$��zk��i�Ĺ��, r���Blm�
j�ttH��vK���q� rE��N�{@��cӒa8��� ՌkFQ�� 0�q��:�	�����7s��N�Ϩ���b��S�d�Ǐ�ū[־�PS�C .�Ȼ{P�i|�8��DϿ�`�@�*���B����B'p��(ۏ@VzvJr���rXu0�#U�W5 tY�g��9�������U`ݻt���S}�����]��4+���Ȥp�:�_� ��L�����ޑ���B]�B

������I3��)Y�Yt�����]ɏ]��]�u�fr��,�w���|�O߈��<į�X�<���R�2��?x���pNE����z��
�P�4	]��>��mZ�Ȕ�}����L3A}��9��qS�D�`��O��g����
dĈ�p����b=KAi>�O��%��!le���xi�O;X��"s��s�����9[R8�SKՈ�FT�>�X8Fń�����2&&&<��˩��m����)6eA��	!�yD�ews�D����9�7��� �=a�'��Y�k�_��?�;̖���3j7SG��}S�G}?8�xX��WH��^��V�b1?|�m�q������'����Ĕ�B͊���{p���t��ԯTn��8*��I�}����(].Ǩ�A"~��Đ���ej��(=��"C3((n�<�����W�9S�M�e�����1���~�)��S�r��'�\}��\N���X��"=�Aq���9��_��n��J@`�@��CZZ��{6}E:q��
��G������u}��?��1��_�v0��P�j��t8��VSS������ 礯��v:T�欭@8��"�W�Ƈ��Y��s�7 �.LZ�MM�I�?~�G��1f,ժ��Oq����҉��D�Hr C0}�իW���s|j�+���,�eao�뾽ZV�
�q?�:���t7	 �� ڢ�� ��:�B�Q�u�~b�7kV�L���z7~N󱢧��VyVo�U��W�J����[���q2�u.�^"x*jZ����W���ª��r��k��>\�[�m������a��9�C��2`��9ن�&�g��2��֫U���q�_�-x4(�r-��_�gzx��蹏��Y6rKGē}�*���OV����u���MXQO���
��<|�]�8XY����?+����333K��I2������`֨<��WZ	L�ȴ�vi�]�����N�Q���Q$�~��;hsp�d/�[d��U�a��	{\��Yk�<���/bh�bw@O,�u�'�����~����m�ˣ�¶;���9Ѻ=�֐[���ζ/�]��+�/�p
k�g���Ө�D�a��v���h�3��D�9�^�� �<�MhN}|[[[7l�[V~��}�2z�s�n��Q쐘<1�m}��@AF�O�mV-��c6��u)`�Pk|��
>��߭J���A{g'�hj��N�[��s�<�.%̔UvS���EN������9=<"'}�B(�$ r֣�����)�i�(]m��A�J��m�����ʡH0˝�åa>B���>a�q>/�Ұ�J���B.�Kn�.M�f���d�+b���)��k|�O,��ciyyfQ��	�v�z_9 u�k��Ћ���D�n��K;�XlA��q}?K@�� KQ��G��|�+)Ͻ����!�Ƕ�D��c���j3o4���_�c/M���BT��]�gj��L��E�n}�2���~�ʂ������c��I*����a&ff�<;m�\\���PJ8.���^ ���б���@�-�Q�x�c���홚pb)~�K�z��\�VD���А�1a�=		���ʬ���Ǐ<*�~��
��y��s�6	�6K"��O�'&9�x \�F�MU�y\<��lW��SHL%���G�����P�!Q�k������@M�y�b��#'u�~���\'Ćv(�"�Ç��S��%E�g�k%#�L����Hvgr�	����O�87U��I#�9I��U�.�ەcX�5u����G��1�ѡn�L��S�F7���YI��c[��ј$���S���Zȣ��e>�,��SJ���ode���&k.�=qUܤL�*���@̖�%=�x���B[甽�օ�\���^��@:�L����0j֠�����e	*���hh9ҟh�s/4�J���z�4w�@�����'E����CD� '�#	������@տ�K�<~aՇ�+[uDL����ys--�ᑑ�I�Y���R�k��}t����h��L�ﺥє����S�(�s��4��Ż-HՒ96G&G��!���d�*d}�`e�`t�E���,��/��[z^:��=��J��}j�Y�yՂ<T���\�En[~(<�&B�V>-:Q�V��gb��m #��v�0��uZ%�h9�aXƘ�R�೻k%Y��e��^S���,��^���MO��سsi��T�4�����jA�9CEDHB)~�j�	�Π��F�ݣS��W�LL�@���9[�I�R<3��w�Ao���C7��ʹ������e%�<$+�F���J�hDC�A�(�)O:�G#�4�&���DscP�K4.R����x��hɄ��-��� �&(��@bdK�㭻'n+�n��gfbb^5��W��C<����Hs7�_�x�׳Cl�ǀMǑɊ��m������7�@�-/���'7�js$�������R�ݚ��l�6�k� ��f���S4�K2G���(��۩�],��UT��������:��_���h�#"��:���WF��� j.mr���!T,�R�Dp9�
;��*�u~�K#?��IQ�$��h���\KP��Qa��^s�V��a�����J����F��T��h<wqQZ�Qua���#��'��Z��WWW2��C�^�o3�-��=�����}m�@���.�Ǯ�����
�Ĳ�?�����x?zQ�M�CՀ��v5~�����&= mP^���~��/���Q�&&�A�X�1~����獚9ny��39j�9<Z�DMǸ8�E��׮hrݞ<W�u�	@I^��3j��y`m���xQ|Sm<G�#��&�ˆy����;��ƠW���,�wڨe��� ����H��o�&_�7py�y'����-Ѯ.1MeT/Y#����:�O�a)��	і�P5�\�&w@�H O�14LMi/�J�S�m��SļԽV&�brP4�&���Jnc륻Qa�E��_��-P�;�4��S5VxÍw����&�f�ϟ[�p� ����(kt���q<ּk�N��-PP��n/�����8-��}�ֿ7�u�86�0���~i��g�{��T�P�'�Ⓚ�A���9N�.%����U粹��UP�u6Q����k<�x�����C�
S�Qhܨ<��3)s�N�,F����gj@��� &(9�.��P�V;"ö��\�my��5A�
\��Y�ʙ�b4_)'�)N��(=�Ͳr&L}����SB��7���1��?�<�u�GM-�u���%���]. #%eCU=O���v�o��j��b kf�?�Vk�>I*�1{W�j��|���i���Z�a��<����B��%M���s��"��
?����vj,L6��
6Ѥ��Vrw3����Y]{hn`�Um<�;�Gu#�ɠu��Y��\8�F���ۏ�*���ɩ�S����|�Ԧ���N�FF�GƘ���kU�2lk/	�Qw_�"&�y��J%O���(����l���&��h��ut�(`'���h�v\-:"���i�/{�Uԯv��Q�`#�7rrrو�%n���X��K���|�]ȟH�p������s�h�����r��p�eP[���Z���&��	B7İ2�9����ke�* �p�Sm���)��yv���s��T8<۩Yz��eZ��� #���%#+;"@[�[�;%����LAT���6�SmJR<�kU	�b�ыss�v��Ҋ���e�5S�ˏ���S�p<����ohƾ"~�Tc�V9��k�b�O��	�5`pC������ӯ���0b����)�k�������᮵�S����q-����lg4�mNh7��
���9���^���LL������|���"�_K����� �"q �(��&�Y�;[юEA�ai{�V�)y��tvSc���`�Oh�(^�  ���nOU�"���G%�y�@.�ɣ&� ���@�̹������3mr�oy�� �l[�^��oAʻ��m�bgǻ����R��TU����Ͳ^�unp�XilCt��4�2��z�`n�2�90��a��/1)�0�
Iګl���iS�3u��l�7��$b2���J��LL[(Y�Y�o0�7֥� ��+Fvp S��#�EG����vK�{& ������WT��_eOOO+k�U���\���n�x��^+Y��On�]����� �x9�n LLLg�_��:����%Zsb&ʹ_��M�?<�;!�ڡ�����l���#�Ȍ: ���Vf��ǭ�e):P�F��S��P�c��5ǔ��i�(�h�R���tT�����ï�,uTU�+��^��� ��(\.�X�>�ӓC}���m ��U�EZ���c�N�Y܅]!A�9�B}dd����x���Y�`\)�������O���.=��({b�}8�%�2�_�@UM ���ר�%a���H��r��x�D)����a2�ȘQ�j��޲��ڳo ���[NԷ������UUU�t��ψKH���M����-������,m�e	Ү��������c,�`儺���-�Q���W2f���/��@�&/��ݞ�L� �%r�������\�������3�c|	���0��[ޣ�O�#�K�.dvﶊ�R8�86C�mh4l_�7J�l��%*]up}:�o��DR1�#�A��}�uƲr�p@��D��o�a4���Ȉo��^PSS�[�^P���Χ��{�N�&�5��M���s╁�$��kW�����P��9����U@ےS�Z�2y��]`���U���|(�����U��	�c",���^��������F{�P�,�ge��7�N����b�qxBa���O�ftۙ~
ٽm���g"���֞>}zv2e��A �
��г������9��wm��r�����vq��mC`l������D���N_H���������0$�~y�Pn�eY�]nt��AM����.%S銹5��m[��y�{i�K�p��c�E�xT����!��� (zg���~r������b�`6.Hr�	�ͷ�Ir�y��,����u�c�N�}��M���>g�o�U@����T���{�T4i���&�T����͹��b��9I^�� s�~B�٭�Y����>��3�vJq�y]g��ڟYtï��u�M�3���lN��m��uޞ'����<t��S�9*��K�	������mDc��X��a�@fҮ�;����!%�f��웥m�j!G��Ͱ\Qu��(�a�/��RVV֩�^x��������ބY��^*��sddd�I@��u�$�seY�B+��S���YV�a��L���l\%D**>�����xiʜ���l�Y;;���P�P쏋.�2<$+��}h2��t�$����U|���ð��pbR�h3��(�X���Owf�|Ny+U�����98���+z$\�Dϩ���l�0\��\u��=	^�h�W��9���͋x_�{��5Њ@�� J��ؑAUwOp��&�L���J!$tXkkk�)A�v�)�#
�"�;�+d����o�W�Jc�AK�]�����oy�׈IgbARp)�\vڟ�z�B+&�Zվ�ë�z��6���jT�3:e�{ssS���P��Aٰ�z���ÇWH?*�'���t��#d��o7j����P8���NVH�*YnRj/V;4,��!�J&	C��hb�s�v��1�g�*�P
'�&?� -.)�b�R��b���o12Y�[R���Y���|ө�3��yy���y��)%%|�7�J��d�L���&HoD����?A1Ǩ�!�`��eb\�{p����	Y(-m!������'�S�j����;9R:������}8�UO.�K�b�?���v��: *�l\��=1Ra��Y6���	tL����X咨�Hg!�DDB�	1]�%#6�̴&����MdY'L-ݯC%�����y����w���4��������Rn4�es��Hm����?d~���-e_'�Ǐ�H���6��lƵ���b��
W��~�u�޾҄� �XwjZ�����'ۤ��Fz�YO����a)�7�惰�L�:1z��u��"M�G!� YP�� '�Y��hV�B/Qx~�W-���BFA1� N�9��l3`�?ˡ�;W�z��I�N�p2[(�R,�G��}o��U�]xt�-s���X�x�.��J߈��ٯƤ��0�E
YW	�19��mk�j�em��as�1�����x�~~~��m���#.�5��ԯ��S7�Jp��v�sxdhC2��c��sJ5�{����.�X-z�I�P>��лߖ�"���b�BT�b�Y��F	N�VH �L�|ѿx!���dB�ExD����lc6�2�̾ք�E�HrAb����qi}i�!��(�����2�Y��/��YH��I�umi5�o�_N�(J�XTTTɥ��#��s��Tzg!e�n-�(�Y�����TPP�/���,�C��i��-��Ŭ��;,�fxH���mS=��D���2`#J����is�8D}n:#�7a-������@�6?�W���U?�O�X\'#)99�X���_5\�u���D�����++�g$���1�p_��;n�h#j!)k3jsڪ,�|�g�@,}���Y����D����f����"�9����y�# �r���hh �{{ۀ>q���XP�:��T����zaw[XX�k������N|�>+�M��~B-$,Lq��=��n�8���/���b�`�`	�m_~ä�x�ڗ�N��
��""����,Uu��$�^�f�]=��߯R��y<�]�E@=�Ĝ�<����-`Yb��8j~���ܱT�pV>����/`�:�2��=��ػ�_�E<	u6b#�C��O������?,D���	(���*7�0z����鵡v�-�>+@?G��~���N�������������o���*�V���Q �:z���̌�w��D�����#��J+u�i��cbff�q���lc���=44�~�u8-�iJ��/�O�d�^]�3&&��k)
���@%pmܝ����?9*��0�fd%v}n������>A�EX�m 2�hlP�BOQZ�W��>*���N�����G��)�
��A��cbX˥��ED�2|/,���6��\��Mr��� /���"�e�L�.�R�� >S��B��RgT�I��!�CA�MǪ������y�� ������t9Zނ"����}}��\xnϱ�pp����O?ݞ
)��O�1_���?^ώ5F�ܞ�NÞ���Ha�N~%��9� � \��,i4Ó�K������M�J���N$	wI��GX4}��[e�aC]�#G%%������۪�L�Rrb�y3bc��r�r���V��[G���,T=v@Ѯ�Tť/�z��V��#�����fเ��a]�Qk�ql\܂F�os�h�Ġ�����*u��6,��%F� ��b����4^�2����E�r��q�����'ۅ3��1�7k鴹�I?䬤�ְ�����D���{l����'���r$�\�-�A��GU��3���4L����� /��_��;::�X%!~��p�������g)��7�qg����s��LDE�X}K����1��1/$pg'�;��HD�ۼ����H�ix�|q��O@)��px{WW���	��o9_ǌc 9�1(Ր�
7���d��j��HyQ�7�<=��q�9[(W��{�����Bt�#D������Į!0�1 dL�M��YrZZ�>'����?p��'�g��i�'?'���G1(�<��#���\�������$<gn�1�N������'V@mw ׽�=^%���;E������),	�e��j�k�b��~:���� T��@@`�/`�ģ�9��xu�AC⇛�$''�%#�S�9ӆ
"Q���������ڑ��2�CF�L��iv�h�5a��҆��@�mw�((v?y	����g\�����ҩ��wc�UHӸ0/�5^1��W���g����V�B؏�ѧQ����hخ�M(h��ֆHy��U��z>��GGBB�{T���t�g80KQQ�0�jX�Ǡ�`���4�cE�+.4�[K3ns�ק���m�>~�_��2�6O����۳����c����x�p���'����U�XB	��6n�Gb�J�#gm<�UVV&-�))Yu���=�!YW������Ԣ�S�f1����zW�͛������5Z d������y�D�~�F�b5���Ѐ��(݉m�d������;���U��8뾄e����>�hC|ZZC@�:����`2�B{-(P�R/M��4��D�qJ���,,r"<:��O_F-; 8�.;i8T��DEY�&G6˖���[`���5*����P}�*yѽ���OK�o���pu�E����wDԅ�hZ�,9999,�" n�����_���6��'+�&V��� 

N�z�28�		���j���K��5�����0=�}�����͜�$�ಞ�j@�f� �Hɜ^.�0���|r �4�芒֢����zyy�!��Ć�� U�U�f1L-p������F�=%?�8��v�;HQ7�ӷr�������*K߭�p��4� f��p"��	^��{�-7f�y�@J]�ޡ���V$����iEh�x�������������D���$"2�=��r$�p����4��H�S�2,�����'-�ИQUU�l�}��ʫ�9Y����ER�~:Z�
u�U w�'�]DD��b���"��0`��0�5���3>ˊ���	�n���P; X��f�벉��s�X��N(���sn���d&���[�Z�y��ĄT��� �F��Dܜ�q�������7��J��Ծ\V�ܴ��0O?��'H�(o�����bwX�Z���a�*m�h҂�o�b���ZܶM󳋜�V=>IK#թu����;J��m5�$����Tm��h�
�H��[����E��kn��N�ONN�.2۽��<iѨ��:���ҟp	�Vơ�8@W�4��l"�0�� ��%���+GJ4M�;�P��]�K���1z���� p�r��{zz��Irߦ�%���z�����:��M�c_&b�Z��HجƘl�K�id	R�;ε��T�aP�}k�Z�ι�HU�9�`���a�-�[, [
�=$�˭��
M�gb��a���+�rQp_� �7���z?C/��9��]�P0�i����<�-,<���]ㇽ���Swo�E/K�c�	��?<�jzZ��>9�h$l������9>@��wF�E��"�?��^Q��ub]�]]�IE�h�Aokk+��/N�z�Ѯ5�U�^%0���z�)>��[�bۗi�1����G������t��a�Zն��o)`MkZ[['�;&����>7A]�qTR��;�;~���< w�6���������Q��M/ r���|��hDQ�f�6&����]���k/���{+��Fܔ�x���R�Ԗ��G@�BT�\�u
0zP�����Iݍߊ�>:*h�i��Nfbb��}�y^.��L�������穓��%P�P�?v��`T�,F i�?sZ���}�_ѳ��G-�����BS�uS��ךR�x꟟-�T��e+�i�s�LL��0ʖ��y��A�a�}`А�b�t�3���(�O_���Qc##bi/tJ�Ĥ6�^��2C1�����^'w}����g������%��x�Ǥ�� ��A���=�}
f����˗/�b�3��cf����?}5�%�^�fؗ���9G�&�obc8��o߾��Y�����@YcZ�7/K�t��!�:img��k�~FFϡ�����M .�6
�iEFFf3�Ɖ$��ȵ܌�~P�Yq?�ێe�������|�U�V|�����t�5}���ۮ���j2��`nY�\H$�k�̠XB/{����W���3��ଯ�'\���RwI���s�&�^�ޜ�>�	���́'d� �6z�bVt���V�ii?��А��na��#mUj0u}��_�~�<�Si�!�����`�5���뎶��\_�B�����8���[N������/k�2�����ϊ��r�M5���ӿ�RI|K�ȍo~@���f�A��F�KBB�ԭ�d��_ݘ�W�p]�Ԭf�R0(��O(ũ���ޱx�>��#�^�ux$��4�b�h���b����J�ۗ	2�!�iל� E���Q�����0<�lt��2�Z��E��ю0RQ�xer{-�dڠ@V�{�"yN��.�+�qqJ㖕c*�J!�N�PB���s�Xv�9Qh�n���� >�>����hUb�~fZ����Q�$,4��o��X}u)F**�:O��ʍ��4y���1 ܳW94�?�q�qZ��j�������KBf� �3rD�}��@0�kV�~0�I�DM��<j)��F8<<���?���.���1� x����*Rͷ7����O@%� �Q9���P�룢����M8��#�s�)y� � �!$���XM�Y�6�51���e��2�0`qII�_�R'��BO49ͰH��UU�A4qHH"�w���edd~Bhy8p�����4p�;��R_q[�t�૙���!��Ͻ�E���������KU/.�����!!�.*{�F�&N�=����"r;��WU]#3#�Y+�]�7�}����=�KJTz}���t�OO��}fO}2(2E�'qQ�$ss�b=
	�/�",���:����}�'�KE
_Bࠛ�[J( $���Qy����=��J�q��N,���*�ά��xy�.w��|S��R�1#dr��u�]IH�m������Bq�]u�]��V��Y=���"$$,��
��²��}��,]!GKpr<�>ܞ/}��=�����ֿ����CW�>/ח��ϣ	�!������\�ܐx�b��f[�(
v��زF,,8��WC;��W�5*u���'跢	�!5,3��9I�(M׹<��������↟<����$J�']!��������[^D'x3k&/�n�����i%�t^S +����]��G*Œ(F�I�Vg���π���e�iE:�5^��^��7����8�˨�ѭ�m�#��3��R�
3�7�ޠv,��l<q�tk����!%�ّ�y��%���[���0g���S/jd>6��y��݃7�`L/Yt�]��-��wŭ|8��a	���9;�n�F���,)=��L��iq��ui�ŋ�����?����x6�������_�QK��onN�cX}�#��%�h�t��m���m�K��T�Eaa��FA�^��/����V�A������ӗ@S�����d���*ɔy�5T�"��d�2��.B�kLH!dJ�d�<�y�K��������׻Z���s�~��|���9�#<�R&�=�/�42�]Q#m��ֆk����z0��Bn�y� �V1�d��÷�f��g#��'\��������)R��q�ƍ�;�7�:}1KNXLT�yS��3d-��o7���[��Rܰ6É�����:���1J؏�V��l������R��<��F�v��LSGdRh���)�����=�X�P����S���c���C�{�2�����hCb�r�ߊ�A��=�Ol�OA�V�[J��#l��Q  qߴzJ��#k����	�v��LKS�g�N�ph5�~������K�����c���R%��m����-�3�cʿ�K�cà���sM�]M�_͚u��:������h���ջR	f�w��&~~쑑�/�ӑw�(�C�/|� &a�jZqk�qj\p��h6�"�GR�GN��p#O��m����:�.���+說�֢"�uB�'O(�6b6�8��_2����$�y=��V���{�|�Y��j��������9��ӂI7)�x�ˍ���g�_L���3���V[[�W�f�>���&!�9�K?G�qsS$1)�\0$on�I
��U��6�4��3�Ju�u9��������>t0|+g|�:��U!�����p�J��5�5�n+��t��/1��K!K*��y��z�PY�_0h�	7���
��=�.�����K��]<PRV\Xxy��<j������tp�Nݎܧ�ϧ}_�^�����>Ur�Y�+ �����f���v>'{7]x�����iZ�3�d!q�P�w]QY�Ɗ|Yľ+6�z�C�������c��݊�2�����w����Π�Ҵr�r�[�C�B-^9y�5��Z�������F�22u���1Q��}+���A0:����ECְ�S02QЗ�tU�����-8S* 0jc@NK��S��t��r��8[R^޼��F_�'\�,��d�R-l�Be	���/n���d�^G��a�ժ��_J�fج<W)4�5s�~�:�3L�b���7���~n���g��)E��[��ȈF�$�9U��xbp�г�Ҵ8�!���&a+4څ(��!�����Y^��󴴮g�2��d��
׽j��5����h�o����Ce�܃�ß;:��/>�\�.�Hi�4,�fE��	H�	���б-�АX��� ͣ�ZOGVB�f�;pB��� Hf�&T$��H�M�[��t�򜂬��La
��]��L��A։$��O<~,<��t�-��-�ZCY���l�<�춴48K���*���KgfZZ|�,V�Ab,&���ꔊ��H�|rہ����������WJ�K���d�s<d�������ٽС+dAIm'�^7r�C�y��>@�վ�Lx///O���������W(�JO�5ae��^��7���L.A�>���v����ZH�`1�;����P�f�h�"��S��i�%�6(my"�Z��b���t���i��R�� ��	q��"���}���m5=���ޫsy޲�_����D���?�,��s�Q�*�p��5rޣƊ��Y�T7)ף|��zn�^�54�E(�#����l���C#�͕9i�-$�PY��=H�	a�˯��Q�v�&%a|�SEN���w�� ȩ�X[��\#�����A�A9:p������[�Md`�P������)����yP&��8��M��L��x~M��\v��~��+�*
[}|#��Z/Y��U	��&���C1f�w�"9�Kᔃ���~f�F�UZZ�\l�H�,�%�w��$q�"�꾉�� ű��d\b��ow��%���,y����킾��XRbi��8�S�1'�*.iü���v����ZP�R2�3�ɈL�v�MK9�P���cv "�X�al��Ȑ����h�H���>�`�����Œ�{�.C碕-^
�0c`ijg_�3��;	�����Ni7vu=�����ӄX� p�^����˵���UG��炻���ѐ���ʑ�a��T@�A��y�e��(�-
K��ө1�w�6/�)O%##s����,~d�|���>��Y�A�Ӏ~\p�lWi�"��E�%'_j�#��;��,*zZ�����<P*���A-jA�3��`R�Ix*i��W����<﫪�aV{����0���ןC���)�.�J��꾀52H�`ς0g�����Kѿ��}}w����A���P�*�")&�l��@ax��)}թ��߸c&��w����k���|Ԯ\�$B�
 ��� ��]� �(���ɉ��������ƵLv�IBP�6U��%:Rv)Z��:R�����'K�lA?��,��m~�Aua»-���͋�m�E����A��̘�.�"9*���Vة ������H^U_��u��GJ����,*�[����\��8�\\ L��A���l�dD�����/l}���\�[���an����||XaX�.]�cF�47 ~��@�?�ԁ<W�y������D�ټ�
)Z�s0a����T��Řb  � ����ս�}`w��.,�lGT��_&'wW?C��Eí��ш&�����	z p�J�m~K����?&qk>|㛉���5Gv-�����H���H���`�^w�/�&i��y����Nj�k�s����1����D�+$�zuۀ0��<�A"���G�k
?�P�9ȹ���C�)���yDb��_�u� �͓�0���;�>o��x�N3
*�t�C���G��g���~�����V��h�����N��CK#��y�bF��{K"ș*S!&�U~<n���ݶ�+����[.�F��cb�}�j�5.�ݶG_��e���"vY�;��9"+��Τ�f�i(��%<$�ur�Ɛ/�������HE+��F�����b�g�gz�G��n������������_Q��@j0����>_^E_��`���zT:��2�HIJ���q��ܭ���?�s�'�L�I4B��cu�6$} OQY��41f:��e�&9�$�����4��'��1�����{����D��R�>�J�k��G�
G�=�!`�*A����1����`����u�B>k5BW�����~�W���� ��<�����+	7�ԅ��;�k�=F�)K
���G�����(D�n6�-��޻�HUݨT���% ����B"ӭ2�[���~5pEe�&%L0�Z���j����+�#���4=�|%�� z:ܚw�żX/�uD��X!Q�B�*�w
�
�m~��Ǖ#��e3&�h"d�zvn.��ӕ��?�Ԩ��
��5�Β��<Fጞ.樗/_N�"X�|�n��s�����p�r�Υ�����zЇ�
;?����5�}l������Gѵ`B㚦~��kt�ʹ�8��ӌF�z2{���~�n�����h�iK�<8@���混��|h���U��M�B;��4����0ԎeС�E����ڝ��-(߿�%*!H���ku����h�ǌ��̠9�����#���)��
�E�N�;s�UJ��9�Ԧ�����[�=�BL�[�ѵ����0�`�n� ��Y����$?�ȸ�'Lο�x��P��>D�]���	���=ZbiJ1-Z
RZ����v��Uf����W������%Y/+��l�����B.�!��?6�����)p����o��$�WI�Y#��;W��o��X�u�Lo`^T��b-ww�$Na�@{SB�=kmmM4�?�`�����$!5x�=��Z[^vy+p����+b�kvnzz�ka�9�6o��}Av{�D�����n�n�k� �b����n��L�-!1!%EN��D7T�8j��/4P�Yz�״���'lɃ �-)&��kO������1��(1��A����X�"#bPr>\������ߗŖ�9����W����&M�L��bL�-���F���öN������Z0Ů&6������9ڠ(T���?
u�(��{�\��*�㹷��l.Ҹ���������k��K�L�o��G��ۑ��е��ފ�U��x*( DbJ{hNNN���H�F��Ɲs+n�-6�;��kյ�v�gϞ9ܔ��OjCZE�-��ۆ�:���(H���f�i�RǷ�7�0�E�8�"����A�@k�����F��ZuSl���.*��N��n�����ǼU&��K���O�C����U��q5O����ȹJ}��x�7��~��*�'���S�>�#Jy<V�T\��g,��weIU�zYXNZ�
	1Qx۹�8�T=�5鶹��a�j�,-�1�1 x\xߘJk�����E)�p��3N-�"�R �'�A�qf�\L��mn˚�
�5�� ƀ5x�A�#�����#/�Ǎ�X��gw����BTw��Ϸ��i<|O�_��o�pa�<��<J����>����/�Y�qe!�Ƴ]�q�H���s~�$��ƕԖy_ `o�a~߂�PJ�������h����-��C�X�6մ�jۗ�/ԅ��fټ�M�|�VD��v11)i#��O�IC��������p�y�}��O�Fc��~�A?�@�����h���M,,Nٞ�?�x�모h=m6hC�<���.J2�~=��E�4U��W���B��#	�dl��t�������_��ʫŰ�_YwFS~�T�p����xʎ���(6O?�e�;0N�JR<Q�	m0����ur{ �>[��}<j*R�dE�x����-P�bok.��pr��y�g�M䝣=%��|�ʴ��ߚ�S*V>���.�����`����*�۳VKKW�	E�h�@�"�;Kк���� ��W$JC�����cv�����n3��tէ��	�[ec��N��^��oŷ����ݛ"����ի�k��+O@�c�(>/����&�}�*���i)y�Bw:�v}`v�����K�D���Ŷ�葦������B�l��b���W~����m�$�ѝ����'g��)8:?��n�i�m�#ˮ��{�	��ĤKf�O��t΍�����P���,>��q�6ԯ��e��s��_�u[��g�ׂ��Tji�P��#�	>�}�:׿�&#p�4���n���<���	����1�}��O�>�����<����83��9��{��o��,:���V�s��cY�@�ٝ^E�R��z�7�O��o�]�Md-�-{-$�P�4?����9t�2Z'w}�!��\���	}�}����ܗ]��`�Z,Ō�7x����u��U焆{S�;���`*�d��޽�&���#��|6��0`���P��kH�A =���U6�e�a��ﾛ���
��g�N����Y�h6n���fC���G�be��D�m��+�f�%�}+�qyIF*ME��{�`u���u.Ļ�Ľ��y@A����*��W��-zBJ�B��9SnѲi��ɲ�S.��%Lx�����t�º���2�];:�ϐ0Z;���K`V��pc�J��Uˎ|[pe�r�[�<ܝ�h�&�n�W��-��Y3RN#�᫪U���iŘ�V6I�e;P��bifO���~�s]�}��%�s�\0,�B8#~:k����"+��R�/md3ML�?��!Ѳ[M���p����<��e�9\��'ʰK2;�g}&G���_�!Z�Ko/C��@��#���*8�k\��^/ ��`�U'����,�� Brʩjҭ�31u����ܱd@�^�_����^���b̔W�1�����
���r��D�1�)�_�:���w���u���X�l�|Od�"�����i/\B3#����м�^\���f�E6A���{W)�xM���#����O����}g�D1��g	���1�t��+�Ɖ�� 	��'��x��L���6MM� �b�	L3�T������[�b�XB{Ԟ�5,n���gx�t0���ߣ��v��P31faqqR\�#/�T�r�n���Jj��~�;�>�͒3S󨗩��8�F&�%�m�B�k�@	 �S,��ڊ� �20�KkJ�/��:��LCI�g�9�Y��k��쑽SWU~_�͒n pF1����z�{iɮ��T����[���Iե�g��[�#{�2�T n���J�!��bV�=�ťw��TUU�$--A���no����|56�+�����2o��RO~�q��!�	[����AʴЈn�/�[s�K�����M|�8h��V��w��E�"�
V��Tj�5����Y^q		-��C!�I���%�\s���*߰��=Z��PÌS����I7��P[��<����0.{0��+^�MZcj(%�4�bXS���;�s�ܷz�(�pи[UEq<�+nMK��.n%�P�*0��±��?��81��xS3~��ɝ��xZ�R�RN.�R,b �c�{�-_AL��k��ڟC?�.�g"�8����3nx4\^�
#�(�)s��cn����yb�s	���&���#��W߽�����:H>C2Ԩ�


%g�c10����\۽�	���C����;��^|���e�X�1/>s!T<p:�%�0�kXkX\P�X�wk�{�tA��h�.��"���'����̐S/�;���,�M�J44d$�m���\�e�C}!k\b�Od�?U鱓�L:U�b��h�l}Ae��;^��GV�!rSS�����E�M@u�m��WإG\�7��P�Rs ��������g��u����7FԢ����9���+�w�ueF�]�� ����t�ҥ?�����.=\nQ$'�I�N����b/�^҂�j4���L�hϻ�V��F_��ᑜ��{�[�HӲ�6�u���G�G��N��BD��?��L�&)|�Wm�:O�̌�i�P� ���Dpj۶Wϣ��v�����)�Y3��ΫPWY<EE0iz�}ѦՔ
o�CX�d#��Y[��[ь���_Wm]>�]=;�	~!����<K����:���kP����*}id�7��#��%&
"eiJR�j���N�p]]]�y걯��! �C���^z�kx�`�T\��2o+B����gMӓf�&!�e��Ԟ"QR]���f"*؍T{�bn��p��l�`��7%��M8�筦T��\PL�g�\�QY���c�e\4d�2��%��J����y�n����w�����ֵ��a��G�'���R8�@`��Y�U3dq�,!�C?ґ�\YBk=m�V�g.[D�{���X�C��O�9/��a�9�ɍ���_#!"$
@6�.�ٚ0-�㥩s�yWt.�yWTd��oؚ�Ԝ��b��򑢥|m\���kkg�ք,'Ǆ/FtJ�S��D�5ł��k����x	fmu�*����x���$X��(P�^'Kz�P����,��'�+D�i��Y����*�p�3y��~P�0�@���q��Ρ΋f�Fu%%��go���:R�C1��w�u[����l�p�Y+W���h�6e`�ڗ�Yݖ�q{��ʩ��')�˗��,5ى1C�2����j1|�v�;�
�)�� �h`�LE��c(h�Z�v��ګk�]��~ةT�!Ǡ�o��|�9�rhi˻��n� �F��E���{��Ab[Ma~��&��*r�f7J-�VB��qݫ����,##-b�;l�M\\^�B��磔j�ni�Q�=�)p�n?�(�
��l8�w���x8���)��T�ST�Q&
ďDH�vx�ܶ/�מ�=B�sA�3�N'���Ҽ�|�b��H���1� ;� �3�'�&���yIO�ڰ�1�6�u}�p�b��&���$�jv�⿭}n`q_�@�TLn�M& ���)K��bd���Jy��!�d��Kx(��s���ysNR�"�:���O!G��s�0ސ4�b�9�_�ܑt����������E
nh�e)F���;��@�=�T>d��phHj�����y'��xJRm���?uj[ ���Γ��J4�[�B���Ş����:��PȽ/��$���r
`������)���b�9�^��~A�fsh�"q�I��cԖD,կZ$vtvf�`�(�Y�����ٛIo�QYn i@Y!�*d߶�`
3��d
��TՄ��e$�ǿ|�N����d�e�~�P��m\	�<�w��.�9��:4��Ǐ��'��y�����D.�8�X�b-�y�|�&����p�ʯϓ��(�!� zb�����,Z�vX���<T�qg�[�A 6�ef�S@@��2���4hrP�~���$<��@O���'߸��[�����ZE��4�Ȍ�9�<�h�l�}��mi������|zq�:���9�F?:���\N�}��݅Nc&2�.%��)S�����{1d��̟_{ �0*�4�׽���� (����~O���n�a�y����C�ޔ�f��'&��������]٣�ο�cc�sB8J.��Ӏ,�LE�-�}�:;;�<��0d���s�^~`�˃b��
�eJ��|���G�#���׃ɭ���X��G��>B�eW�3P���L�w���k�(��K�w.n4j �Z5�>��-���F�i�3)(����$Jظo�À\����VGG�L�OX��F�bՏw-�4~惠��~�L[����SBH@U��Cw��N!��Pz�������.�sD�͟?խ�\�[�t(q0q����+-i[6 ��>y��h/4,�R������Z��-��+F�% ���*%��݅|���O�UN'4e7H����2 ����$#����j�?���R��\t�ߴ��/�B-���>@�P3(5VYn��Qk���Z����;�B{߂�^�,;cE"���9��^d�����pt{k�YQ��Bs'k��[9��?ڈ� �/+��p�|�4�/�u[l����s48޺�� 5�nB�*"Y#��nX8{٬cA>ˡ�<�-��
���|+�%ed��\T;���L)TiF�˗`L���\���N�|���W�L���B�躴�����7U��3����!Yȵ���V$"��$���(e����(�����E&���F�ȼ���J�Jޚ|��dO"}K����Xihh|4+��s���Ы���������9U�i�����������pJ�9�'�� '`x����#�ED���m��Մ�$�_Y�5�YX��v�	فʠf�aº��}�p����9�R����^mv��imx�&k���}n�91�>����6/[��2��ӧw��x j���U�YfH�Z�Yn]:`٣[��8��t�,*j%�dʨ�h�{=���n2�J`�CB	��NAD����
�˯�����#m�ޘ��,ʊS����n.,/���Ȝ�y�"���F��t��`���i�2���$�� ���U�_�X$���1q<��6-��A��{=---;l+6Eo
��P��t�o�s�i�d�$gӥ�%�yߧ����T���B�p4rRU�����Y'�-����6�ͫ�zzzP������r�_�z�%��]�G�&j����s��3���pcp`�(P��D�XE����1S�d';���<t��4*ZKN��;µ����.�%�)��җ_���.��t*:>��![T��R��T�H�su��`�򞓪dw7 x~ʃ�������B��Q";8E��^F���G^�pf�ٕ4]�������(�#J���к�T�]��8+��9q�k_G�5�۲��b�d��F�9p ��\CS�ɸ�����H4
H����yȼ,�`!l��ۚ/�F�q��<�+�=�6W��Ľl��J�%B%�R�}���]§R��=������#G�qT~��f�RY�Ã��ș
fN��j�0̓��`�ُ�v�AN5�~MM�h���[�mi����:j5����H��u�1e�I�3�;���t2\����bɐ?�c*�9�
Nwg̝�eٰ�����s�|D˦��ּ��-���6�	��_O	�H�g�,�>���"��b��2��vB�a~����\rFG�������mn�KŴ4�<t���T�O �L`K7p�X��bZ���������u�
1�a������b?d�WTT<o���:UkX��\�G��!�W�F)��f��R"d�	�Q���([P:��s��a�A��?�c�}�ռ�x���`H ������K�ʲ!:-L]ީ=O��j%_P�y��k�8�ªrpXl(���C��u�Z���ML���xTv�׀�& ��ƌ~��� _=�Bߗ�:M��`EV�X�P(f����׷e��b5��g���^�,7x>C��nGt����7S���s�����;|�˘YX��ȃ���!�D�:��[�� �@��K�x� Ct�-���$Ci�Kg*?Ѓ1�W������&Rx/��ϣRڍ���,��u
ns�w��|pɳ.�X(�Ug���G ���v�I��65#����F8==M�|h� � �e|1?hap�M�W�4�WL��
��6��v���H22�6X�<S\+�ٳgA>�G�iե��_�+#���� �ʯ��T���Q0�T��K WWkwW�r�Pէ��uO�J@�+r��|?^�	9��1`�����7��BtCg}գz�î�d�WM9����-����/s0��M���l �Ƀ��qo4'M�?tВ�Ǡѯq '��s?����H���!�f����ɥ�
S^��s��8	�]�U�5>j)��	���U�M{��� �L׊ܫD����
u��S�3�t��X�g��F�����v�iOg��.H5	��k�]����Ǉ�Fa��`�UUR0`��E\i2���  u��!`8��w�츩�#U��O�y�_s��w؛M�2A)8�}���:᝝����8m���J���:@�����'űf�-y�hT������Aw��V�ŕ;@�+���3)�֤?�gP�Dş� j�%)]13c�˔����0���L�C����v���@�./4A���\�tG��l��N&��T�,
S���Q�0�ɞ�C�)�/��{8�@�,�ݏ�C�o�!l�;�!�����N[��O^K�չ(���pO�Xk5�	���N�p��I��)�N��#�c@I����ȴl(1&2��~�3��MT�"rH�b�:cZ��
���ب�G��^�~��`\ 
����L@>���V@P�B�:����>M�<(��;�L]5��=\�V���!!!ܮ�Ԥ�MǨ� I�h����Yaaa����*,��Zp3k������e��E�*�!G��ឫ���l8N2�#��;L�����g����U� )z�� w[�,����(&������a��z͑W�+++�ň��L��􇹔?�
	W�0	�)Q�b��Tqq���:0|�/k��?LE綐���K��ZlX��1����Ga���?�H<!�b��'N��V|��K3�?��h5@��hw��-�?ձC��Fs'�=~���Ϻ|�aN�@[��̏T@�s����� p<ܡ�9�����P�b������Ky������\�s3�'�}ǸlYR5{�P�H��i�*�9�{��$o��)ԪLh3�q�+|>I]­�$k<<m� ��4�v�ٮے�^����w@>������ ���ڈ�}��-G5��n���t��k��G(V\B�&�w	M����i����%(��nnnz�ǩ����th9�2��=�1�������C� �r%��,;�t��qWk1f�ݢ�.#6�i�ݼ�?|���pU�i����J�o�/_� Ou-�#�?8�n��A����X�j�YO\\��j���`�l���"q<J4$psR���:Z�)�U�뵡ؽ�,��zz��2�x+�t:�����)��������N3u��6���qF���� J�s;���?�Օ�.*�s��Y0b��Y�X�9(;W�BXcX��W�M� S� ?���{km_+�L,��o���·��z;,6�Kxo�+�ʽ_qh1|[Mc�}M]|-3�C��x�����w�:�,��ٸ�nLZ�>F�3 9���BY���0E�2Q�B��{���~[�{�h3Cڍ���t.��\\$�ce]�b	��mP�O��ﭞI��J�}dgo��ҡE���Y��S���-vX���_GZK)�h���V��G�񮒸G@���-��A�r�>}�*���H����sk�-<+/�Vv�ǹ� �$-~��Czi����e�����[�c�n��_M�j�?K�Ji�XC���&'x�\����d����~r��ꐡ��73�|	��	�w�V��W��-����!M���t?%�2����vs�}�D9�r}A��Nn*&K�b�}*�2�,U���6�
�r��֡sD˴w����VӠf�@hC���YTz`,k�L;H�Ǘ��w�z���P�¥w��<�>�+3�ީ��R	��vvȩ�0���S{�BMpf����������8��n5�������J����p%������9?�ك�/���Y�z�{��Gj�݊BL��ee2�{�W�%������黖��>� �z_Q�6�
ޗ��e�
:x&*��Td�����>>��I=�����}�ɹ��]��ι�� W��m����V�-eUU��h�1d���Y��NN������2ҡK��i^���hKR�5Q̡ՠ���^ZFN!����S�z�9�n���f9��d�ni?�Q4��W�KS�c>������Hb�\�&���D��۲�;PB��s��N�����di5����Եw|������^?Yi4z>2>���Կ�.\��o�#���	8U�J_I���� �
�����{g��@�G��5B�T��%���
��f2�m�ۓ&Q���鱫��f��y���7R
��8LK��|�C��~v2��B�%���!# :I#��;�I����Ԥ�G�ɂ���v�Fc;��t0��}?p���a3�n`�.��F����kj���Ύ�wr{`��8i&+>q9���n���?LuƐ4�4�IVR��Y�Wy��Xh��KH6�߷���fg�Fi�t\��Oo����DN�Ȱ��|��� ���Z+�$ɺ8q����D�௼$SWL��]t(Rp��� +��z@%��\>�8)�ռ�r��C?�⿖hVn�S��*��"����[i-�L�ּ�x񷗜�ж� �6}�����D0�у�G���Y�=C$��8�*
ep�\���e�gh�����5Ըu�DY��L�����)��2S�p���_�z�-�BX�ۙ/ᮻ,�x�PY��l�~z�&�KzW�u�~QbL[��͌)��ז��^�p/�=a����ϡ@t���iXt��I�Ze�<>�b+>RW�?��B�Ŗ�[dT�>������k��P�"�h�d�ʮ}A@{_�],ip��a�񛴗���ؾ�8E0�ٸY�����!k����3�c�òY�����FFF>:N��b�?.�ڣ(��xì��|.Ls8�fz�4��-݀���	Kʥ�!۳�E�7���������������H�5�ʇl���Ż��#�b�R���iH�_���b.r��br�Qp=���8�A�[����8�BS��b��c�d�U�Aֵ
�p���'��?Ys`�"=��(,'7V��2����s�����M��e��k|~$��I
�ahi�כWj]��3�l���AQ�ۣ�s�rf�����e�=�d��nax�,�zsGGG��X{�:@/��[�Tr�8۰x��G��km���Ek%�)f����mƧO���I�����_�#�� U�$��/@Vv,�a:�S���]�v���/&�����柘�ҤUђ+3,@V��y�q5OV��]��R�lȶ�y�w̦���n"��
XU�%V:�w�0d���=��Pk.2LZ��G��a�E�Ӻ>7^�֐�r��x`ds�����2z!���q�x/��Zzq��uu5���FK*�;��6	7N��9��/��7]����k�|t���_�G����c'H�WXxY:�� �9ӕ�t=NHT�,_�w����=>u�ve!t�$���L�$k0��5�F�s�W�BT�
�	�dIy���&��	@;�Voҍ�8/��>��ُ��<��֔'���F&��0���Ofw���,h�{Yn1(� ѫ�i�{=p.��*=�{�ɥ�R8�{>�"f�%��b,�C�{	��y�Ω�]ܞ��ϟt &��-A]bU�S?
OZ�3��84?:���ΨW2H`�p��R��mE}�=���ؽ���n��� �kk�<d;��=T�i����.��c��/[���W��`|��[��<����>^:��öL�a�e���.W �S��>��\ԟ�:����A��ׯ_'�v�o�v�^�#Ij;Q?1���!o|��6���
���GX��b\���0�����ŀW�j��o2�fq�c��+ip��K#����S�!p�#�6���G{q�f]�dI���I ����cs�
H����?��q@dz��9<J��_�K�0�b�`I������B'@� �]�q�?�{��|!�e�iIQ��|���Egk��[�7"�|��K⢌����Y�1�ʺ:���NU�?�u�.; "�	L��z�Ox<g�E]!!"��o��(��TTV҆�'�jh�R�z� %�5�K����q�ffm_{��������s�U���3]>`(�[��/ba��m3'ͬl�J���Wf֖�"岄�<��d]�
���gh@�ܬTM3NV���TWF*�,�gI�~�R��6HN�yP��F��s[�C��(��z�5cF>��w�v���k*�'-�3NR����>RݧȂ$r���[on��U���/�}��YÌ�Ƭ ��jv��������e>O����������2>���;of*�S�u������X[��p�����\�[��K�pO� �V��3�$ ��܏p�u�$p�������ȓ��r'��[s����S�:1�w�u��]���'ud�f���8��މ#o�m�V7�?�I�3..G�v���9}f��}���gׄ�s��jb���BC�Y<-w(����翍���˖�2�ӱ�ı3z���+��#��UU� Rfo���z��]�
�|�<���~8�֥�z�t�H�^N����MX��m��"���2�R�1a�}�V;����7Z��"]��P)))�55,�cZMM���U��N�>~f\�/a7:uP�r���ypo����jm(���^^ެ4��_+��QQ�3m�\e�I������:�8}9<�}��A�%��"|x��h�`a�fNN����i��L[������75Ȼ������S�Lb8��;ZZZNu<~:5�8���y�����77E�9sW�c�jxhGnZ����ж�.t�m��|�tȶez`s�C�J�����hm]]ݬ4r��]_SSt\k��z�Dqqq�Ǐ��쌌��??����7��~k�U���#y#e�R_���/	7r�?��:;;�VT�޹sGDL�aS#�?��@/��9t�E�Ћ燆���
��u"�5s{�%#�R���Iź-�?��V�ă�J�ȳ!L&&�����ٱccc�-H'e�}�toe�~~�^ѷ�EuQ��K��q2��ے����Ui����HH0�Ş=���<9}��g�9�_��`�?��H�j�Ib��h����P��y`a���p³�##�		g����#Cz�i�mőO�ǢQ��x݂�E?mŕ��}~��×Īt��kC?z���IQ�wyw��?����%6E.��%_������ޥ��֯_C�:�R�46*]8YZ[���w|b"ɩJ ̝(���$]�}�wAXɸ�i�Љ��\��y�*5�GQ�v'�<(h-MB���F�B�W�rnp� �({�dl�e�7�����1fU�I"���/)()��>y>��2�_�lW�_��@�Q�F���7��m{{^-�Q@��::0�D�+��_?����k'w�S�o��z���x@�~wljjr�ݜ�1'�8������j��e����ʊ<V��z�<30W�#�$���h�޺Ep�A��������k�bw� 2���R\��\��R�]�O�A{{Mv9�׬I�s2������;� �g�
rI��^�ss3��$s����˜��/W9N�ee@�O�� ��[�2M��g]>�������d�QC��[?@^Lݲ�2_�`3��p�����^�/n<_�FqA�m�㆗>o�"�Q9����%W ��Q�^^��i.��k�	!!'^�d.�v����Fұ��NMMES�CK�SO-嫟�UwX���!�s~�/�h�J�1�F	ǟ����U���ϽwV�iu�:��S��[�;�"")9訿�W �H�͚��:�y�&[1ݩsll3��^:���CM�e��]]�+����w�n�.!#�
����K���Q��~��e=8��h��C*�b�֞"A,�Q
����e6����+KKKlŹ=*��cЉ\^�z�r{\V��gf�<|x'������꯮�pρ��=��7*>���gj�}�����G�˾���Y]�!��^��w�w�!���ӣ�I�S�pop�iFRX;_���MWJ��a�2���
<������³�:ϧ���F�������L2u�������u%%\���/�fh,���?2}qppx��&�n�S_��h��SY�sk��0T�L��A�Ȥ�����*�;��ME.?Z�7,q�>�hFs�s@n�&�u���Wc�IMz)���e@���L8��	�3����j�dK_�	­�����@2�#��%=yr&Jb|������۫c5|Pj��'GY[<+�S/f���7�3�4{L��6�N<��z����,+^�Ko���ё_�����Q� re}�����0!��:ϋ��D���@�y���-�NN~~�ci_�_�uU�ΐ�د�l���nn+1f��J���>[�ܖ��,s���F�ߕ�o��{�4�Pk���bV� 99��c��3����m,45)'��'����A�;���󜜜�Y�����_��6���y�;�e��n/�{�ˁk����y��4s�����a�A�,ZM��n���[��T]·Ƅ�D�
�@r�*�����|ƲY�9���8L[�����ŉj1�%l�Y}֭�?_��/��ng��]�����$�;��1w��᫭s[��������yȚ�(�th�8Ă������������Z\�ZB$�������[y���W=;�$�P�L�T� �liyy�����' qk��ш�ẵ��L\�,AV\��LN`����wK�@P���.�J�O�v�.�ꢹKK���;]�T�H�pC�lbr�ܣ����A�ҶcU],O�8�����M����A`�{GPMῄ˗/�����v5�rY��홗*�躙�3?��`�k��=��Q�4�Rk�Ŧ���\�jH�,�J&T|_W'����p��*���w�޽��u�I������`\����_-Ńe"�W�a^vy��3�0�� �D��"���F��-��5�_���))�Ct&UE���!�T�W�HSsȿ�e������ɓ�-�o����a�����_��6�611���4yH��P!�/Z��������=��&�د4��ś_Y��Y�%��A��&w����ݕ��_�����T���V	z��拊|���@��sl3�C ܳ�I-f%��1�!������w֜}�	��Wz��֠���<04|��bv� ��
������k	y�.����}��U���%Pѩ�1�7s��;�����*苫����˝&�� ��������",F�a=��x���!B�Y�E��_����_x��e��v�/��^l�z�l=8Ftim-	��-�����/q8H8�1aII~H���ޏ�n�Ծ����w�S����FHfKvQ�(d�̲�h��X��!$d��8!d�c��� !J8v��w�ޟ��?=�s���^�9��>���6��{��δ8�:$@��G��o�l[�C�8�W~ծ�U�.�2�l<�R[{����T	�yX�����67@�@Y:::��p[�Zj#��6~JP�r�&&J4A�L��y߳ ՚�(yT�[�kF1ryp�UP���g�[+��nP�~�%@����v����绅�m���t���m���p��h����M^0E�Ü1�j**��`��?��x5����۟���"逽�N�!�w$%y�\�m����gAk�_Q =-�)�[���k�\�ZVޛ)�o%U
�>`0.��=���򧠠� t}3�7ۯ90�M�g��}���T�^~�(��`Feo���Q�ci;n����f�v�8��(��O���&8���^*~6'�F_��* �vJ~���7�z�� �/PL��Ê��Pz^��LK����urdW|���h�xSԛ"ͭ<C�w&�`c�xM�ΝDDD 'E=̍�-[Y|绺�{	�O�-�P,��+��Uy). � .&i�S���~׌�Y{�X��]��ln�115Ս�u�����Հ�@$WGoW�)P�����@&dX����i9�%��oӨ
��Ԃ����GF�H�R��S�����M��Ӗ�V�>7��H��O����?@6xqۯY��E�uss3\�^ a��Kj�s�0&V�H�юͦ6]oڼ8w���i��*|&��K+��ՌNL�M'>^#88�L�y			|s
3+555�X�b�ȰM h�R_�2�$�I�He�}�p�~BV����M���U�;��@�}S����`7*7[8	\VYy�f.0i�3�6����q"�.�~;�&j�a�?�$\k�9�<�.�,;Z)$?E��"�ִWUc��嬚۝&H����|K�u��p�yQ0���k�Tuq�����Ox{����d낍�ֽ�	�l�Io?'�WT9�)3��h#� ��r�`�
��[[5���=�t{�թ��٪�5�l�B.Ϻ�%�W�4$�ӯ!��� 	�Rc�0R$����EL6�U�5�3�����dz��ѣG0C��� �{�U,��7��Y7����Ћ��D�4�[�{�2�譳�=P{\���w���K����2C@@\RRR7�)�?e�<�v��h��lAM�z,9%%%nD"���`�W����,[�#.���8U�0`P�l��
���U���� W���c��g�_�<�h��S���/ook;��Ϯ�uZ�:X��G�QO�� kĆ)��0���-�=�2.���&%�a���G{��o��p����������N`���D6��HQ:��l@�:�����z�:e�=�A�0���7������yM��?��J�Xĳ�J�9 u"��	
��%��fZj`V��_:�J3wf/lؓ��A�M��^�y
�m���I�5$�؃P����W�N�a�Y3r!�.��0cVVW�~�z�n&����r̷6�xUUU8���pf�If�k�U�,����o:��6$�NNNē�"���j?~�1���|��=�l��/�<Y��=*Tx�l������|m���C��xS^J���/"�\�;��7�G(N��o��cggG�������- M/��rop�5��9����r��%|��I%�<+ӫ�E�	~�����	`d�����_��wfgR��O����!cE�7a��\����tڔ��ǗVꦨ<�~�d��askWAGo� �VS�lΤ���TOT>�c���Z���� ��@7��ѿ;l�����
��?��d�76̪i�n�~L�^�Bc[��1�[����SSS�
�{<A��]_F���&a%Bl��=[���ՠ��ԮuPP�uf��&�vx/a)n��"��"�x��a�]������@|�H�Ȓ��%}�wg9��ٙ����	z�҄Rn�kk� �	�m %�����[Jm�W[���ٹ���>f��,��� �k+���@��<��bSw�9�V�Hv��l���E3�`������N�5��L���[������+���h���J��v��_+T�G^���eN��p�����P���"��+`Sj� a�="��W�Ԫ���͖r��[�P7�:,��Uaz���F0�e~D�~��^��j�W��K�Ė*��п��/��h0��N����� �.Ԇ!���mnn�eeRx����L��|˿y1��6�hV<�h,��_qx�zz��=����r��Ƴ��
:i�-�7�E�?~$�Z �GIEE��('-��d�̇���͉?/��XN W���챱�6"�m��9{_9{cl��5=����s��VB�����}��|������t��k��W{㣣���'���Dl�1�߽ �۟�O��
�n������`��2;2ΰ�?����y�_JW�ϩ)�kos޾A	�v��E X��;�;��� ��?3�����/�$8��^���d��7��+�����(/Wo03��#r��d?�h���"Ӳ�/�Ե��C�r�&��\of�2j�WHJ��� B)��$�s^g���pE�ݭ�㆜C	G���tp�Ys_�p��B �%��`����I�ִ�ފ1PfdeQ�9A����V��R�$�|#�Cs�b�~�s��h�r���Ӄ
v_\?(<CD�m`)i���@�w�����5m�GJ򃁓��|�6+���Msء�fX��=Kg�s��:@��F������ xIZ̿�<trq����R22��;��W�Zx
�7q�q6 ���}����::����924ϜK�ŧn���1ZO螵��Q�/���^^�������t�,�^~&s��G�`�c2�$%:s��]��UV^Z���lR���<eX ަ	�WU5W�Œ:�L�rr@j��jB ���TX�EDD�]_��3��fE�C�q<�`�o�GY ������E�6��+u�6���݁���Z�m����	�bN�E�P�.�;.���v֣P頣����Wi/�f+4�D�/7o�Z_���>�Å W��l*J'�$V�b�p�0ο�� ��[s�
��b}}cxW~����H9��Ӯ���G��'� =oo��R?KeOKM%��+,{����Ž��FP
Etx�CYY���*QP��/`�~�T���`�C�jС�0�
&�;�Z�t�_u]�ԵvԷ���k��f�ɬ`��"��^�Yjo�,�*Eί߽s��~�x�Դ�{oi�6���$��bbb��Bv c�e�K�'�l�{x7���~Ω��4��5��Z�f�4��F �ollmk��7�G�<����S����������c��
���g_^&?7[��ק"�-ݯG��X�hP-N� ��:��a�;�k�Og�����ߎ�M�����--�g�K�X��1�ҐAX䛗/��Z<���\���Ѷc�W@�9��J!6�'��G������R�I�` 7Mb������+<f��vBL����L�aE%����
Bəb.<:����V�e�W{�b�=Un/u��邋�q��w
���?77��M"�@��4�Ʌ�ů�E<��c�c ���ｽ���9���$_8t�5��T���ĩ������$�?r��H�W�9�d���SْN���閛5Ύ�]��GsZ�������������	�Ȕ1y��唹x��Б�D<���C��N��A��,5�-�j�u�o	E�**W��]{
�����6I�Pp	'�,:هAm|u��Ç� �h}�5�II�w� �<�T�9(((�Xj=YJhnQGp��zh��6�t��Ф�֋����g[<)/���#��!y3 8�3��O,.�d����U�������;z��4�u?�;�vJl�Nm�����ӧ��`W�K6䇳��me�*a���� 6a���)d�����Ibqsu�I���H��'? 7B�}��ϊ�4L�T�TIZd�aia���e_�0CXxh����L�j�B���QZs^�[�~�qC���r?B]`p�t#kc�~�
:^�<Eט���`ychdThXʍ����\C��3, �3�߾�����KKI�F<�RP�wR�L��Q|~�Ҿ7õ����*Hh�L ��Μ�����*�-W7�?2�-�;h��_���T��zF�A#�4{�vd�v���F�`��A���g���D�3�S$��Hp�R��z���7��o ����=10@;���,9�86�Z]E�	+&����б����Mh	�4N�� I%sS%�v?`j�/[G[��W4ʔ#�<�'��䫄��SFFF��P1S�Ǐ��2�^z�H��1��um;;� ]�JF�a|��n�x���,5`3s����Meiiɔ�!)	�+��t9P����0w�) 4p:���#�
F������K�T���+g(���O��������A5�D!/
��ȟ�S]�u�XN�F�����ݻóc����B��kk� ������B�.7��	�Z-r-h��Bb��S6��p��!�� �M����@!��6���G�<�,���:� ��_��'�抖��A�)���G8E=A�N��4�{җs��UL����- �j��"���}�ܬ�g��:�����D����y(������$����̎z���~����O)߼�}S�{��z��!V%]0Z�hs�i`�+�)��D)6y��]�nja,
�L�F����������k�SS�Ҟ\Y�i &�� ʗeӔ���g+�'����SW_��n\�ʺ�ݻW�/~jh�l���Ҟ^�q���t¼l���-Py��@���O��1���>Tbs>e51�;������/�L��9��/^�PL���w������x{�:��0��lo{�����8!���ɱ�e�p���G���J�@�,�%ܪ���0-34����L�޹�ސx'E���_jWZ@;�b�Z��9|�1�xk�(����h&P�O6-?}�D�y�,6ut��ݟ~z����_Մs����ڸ�0o����ԮmTnv�	�	oa"�!(�?�����td�
���+�����6��iC|Q�S���b-��"JJ�|lr��1�s�VV:�j����v(�S��A�U|<�Q����@���YwQ11��!���kތ�����}�+&�6�wc��_��C�zm��/�xtT�a
�W4�E>��vv֒��4�ge�~�B{��4A�I��IzUTB�����/�6����+	��h�/���U�#�Vl/���#�eK�����' %���v���a�S��'���'3��%Ϙ�����&H��S)���·��c�C�{�}�7^ҭ���44ܟ�}*���ښJUQ����i---q#�;;V��R_�	 WY�M9{�y��XZ���,A��=����r4+�*���:[kb�%����m~C.�O--�)��WcL1�������;;�]R��  ���CCC� �{���]�cKx�����b�"�Ԕd���x,٩kŭ���b{�-���na�Q&L�x�r6A���PH*�@��U�l>>��j/oęUg*X���Ǜ]�uS0��qc213[�Ә������n�Y��2�����+�����!(�D��sz:�}���<''' %����rE@� }ZZ���P'o%UZ΋_�c�k����o��|�`�J/	�9�~�z���_ K5긴��BӲ`�o��֧��l���2'��?����M�T[bz0�i���D�xi��C(�3)d�,p��f�?�׫�����=���g�(�[��>z�S�2�ae,���IPs��m�&
��������2����er�
V&&.�\B�qX^��1]n�PcN< n~,�['�k'��5����_�����'�T P����#�>i�a����W�@���08>25���A��V;d$&�s�IxTxb�iH���QQ�w0�_�Q�ˋ�XXXh{	?h����>=�׮�Z �Gc}������vP�G�W����6\>���F{��k�6}�S�C��@�~���5��k���PLu D���7zȞ Q�^l�I0����:��s(f��s�����0����|t��������R��ɖ�S��
�0#g��gP��>֡^�XW��kS=���Q0��:����G.x`}>���(�n''���Z�q���w�wc�;Q%e159�
ڊƖ��?88���R�(7-s�]��õݱ�5  �@,�ák<f�cɕ�c���x�!����6q�1��'�=���gjurw�M�|�>qp i[��*�i������~�vd"�+gm��x��8emK�@��=�rc>u�LJ��_����Z����PH�k��V��y��ٰ�I1�b�v��{�⇞�@MT@}�����[ls��.��,���#m�'�{�꽈��-��u�����B�eO$��t�rS�����%���r��5PC���s�O51�m"/����7���[���D^Ŝ�mlE��@�B�^�A����N�nh�{f���=�K�B�0YY�_ ?]ٜu5 ��FGɞ��E�1��`���J�?�Z����?l$5<�sm�~T�̢�(��e��A2� ��.�]]�ͦO�۸�>z$\�fV�Mw)w7��ԭJ

,� GQQ��m ��c!�$m�[���c��{�Y����<�;g�o���A�ׂO��(�)��m\��4�#�e-v�G������4�$Z��AQՠ��V2����E�III��,����������������2�9%�~:c��{�hg�U@]��!�B�%/��'E�fG�ONZ<� 5�d��]B�o�k��i����7� _~QN����/����I�����P�����ӣ���D3C9%��]�=v��}B�_Gw�f/tLS$r�����4"�t�A�a�.9�{h'��pi$})���)H�XDZ��ZH_C�|��^��[?~|=�>/S�����Z$�F���˄�u5Yo�vT��у.6 }0����ɥ��7�&��I����.�"���"&�'Jl7���J�B��&��c157��R��6�/�U��ׯ_Bei�*JA�l���[��: �j��N"ZA��s$1W���^�B�3mRҔ��m��՞Br��~ ��&���?攟���s�m!o�S� ~K�4�n�{��n��HY�iik;d�נ��l��̬���+> ���rz��GT:��;y{U��=�o��f�|l���9��O����ަ�#� ��!�2���pQts����1�������U�Q�O�.��>I����H��'�ַލA������e��"�46ሁ�؅!�lx?~12��8C���bAT�����q	+��9y����N�W��@�Xs���	�T���t��J)ƺ��g�������>���W�Ƒ�!�o`�G��g�.ːB�L�}k���*��?�X����EYԋ�n[~��1۰�h�.7PmX�@4u��=z$-A�T���C8D	$��=��-��"�'l'�F5nMo|�>���q%�(���󥄠yT�����cA���m��5q3j S�T�n���ff�m�Q��򝹘W��BB�����Q��N6�
����o���o�(�-5�77��E�V�m�ԋ	�Aí'��2޵�?a�}qv���IDR�,�q�=�D��g�=�	���p�IT#�1���x �Pӆ�G��}���?S}�QL#SS��VB�e��%��A��'��!0��b����v"�֫"�E�76����^I0�����m�?�>�M<�A��~�,'%��LM�v"ۦ���Σk_�}l�ѹy*���7�6��&'2 T��}_Z����.Q�&1�&uZ������Z�:�Sp)w���u���9�����ř��[Jl
��_���_W��MJi4��JoDp܅ �&��`d�|�mZ�\s�P/Nӥ��^�`�ڟ���Bd�xoA�SqJjj�*qI����h��Yw�۷s��*Fjy�d�70�d]����U��mCx�8�<�YXԯ_������*�w�����B�O�e����a -Sޣ�ޜ�4���:���Eg�.>@��߶�����e�p�F�� `uM��H��FRV6մ��:z	�$�<�"�[�&�v,�������/��vA ^���%��]��#{B� C�S`�?gH�ڟgsߗ>���.yn ҅
��P̛نwo�@��),��;]��z���b�T]���#Ҁ���I�]:��c����(�=�����}~�:�_��f>"��J�̍�o}G89!}E�/

؁�;��L�!|�W�ey���5љ�H�NϮX?�8"h���"@�@��A/��WVV�@ �_C���~�����в�����3���4 ��������l�Hqo�v��8��>)�o�����W��1:�g�}Ey%Y����7�P6�VO(�Dj��q�ߞ�	���&���˗�gv�D���ֶ���g��qpp�}zU��L2���ͦ�6��-m�G(��~�����~��A���`~6K��`�"(k�������su �Ն��]�<)���`����p���v�ov����a��1� lf0�1�T���Ǫ����o=:���Xm������`/�}�1�:��J��$	kck�������?A��ihG)=��L-k�r1�I	'''q#�S�/�!��/^�LP�¬��e�z�@���o������^W)�7�i�WH_�wZ�n�H�����ꌉZ����x�0Ѻ��Q�g������G�_	H�J��#�:Z���I�5�%���"mռ�ĳ���Qو�C S�S�ӕ='�L�>�=(<���X��j�Oqt�8J��\j����·�	p����;��
\$@�K��V�d�	K�S�#������v�>��F7��!)"��������O�]I�G�o2�0�8vN���ǵ{��u���쟋dsl]^Y�wS���p��v��S33:Vknm��#�{?���1#��i�>ϜaƉ.Ԕ��'��s~UՄ�-1�A��t+A�n�H����mR�ĊnY��L������i�	vF�J���/�G��N�x��mф�Qv�)?ȱܸ۪�i_�ܛǸ�#2@����.�@�� Y����	[�������t�a�m홨��%��a�μ����!�T��9W�	E^E�P.J"���Mf���ꕊ	(9���� �a�=��ZW�����n��=`���hDչ�Ǭhs�� ����$�b�����r ����ف��� h�k��� ,I��3"����*BC|��:�^;O~���]��e��5��Tk�e�}������f�0�.�S.A�uIt���nxS�V�_w�������.'�I*��H���	�%$�DHuў���pa?|f�VR4Y���B�A�~uc��19�2~7���y�ߺ��!m��L����*x#�����EIz���ʊ}l��9yDt��i>`�R+�55x�=o/7�NQ"��fΕi��cx��~��Hp�C-������b����]�P�p`s�a��h$"������������\����pH��]w)�DS�o��g���1��J=��-~g0������+�-��\���U���	�^;yG3uS/�D���<'!zi|^sr��DG6'�J��9-�Өu��7�.d(��w:}��+'�Q���hiF��(��i0���+-Eu.����k��i����0I%q�����v������y`=p�f���ڱ�M�k��v��y��s)zG�@8��� ��M}�������ئ�͵�MրS������$Y���wD>�M%""
�]^uu�������X�YaW���c��d�`&p��(���omPV�e���l���O>F��nxQ�h��x��p�j �x��*v �9��ĳFH'�vFw0f	xQ`�:of�Q*����q�+�,����g��i³{�v��ETQkӃ.]j�85@]`fw����p>��ۏ��!��m#��!��l��	^���w/����P7)�q�衈8Z�R�9loni��	����F ͫ����hSX����7U�A+lB�O��]��E	����"� [�	$w���x�Z���BK��Z@Q��IF���a�>Ԫ�e��eP<Q�1s�w8{��Ĥd���a���2 ����/��%���gQ=�����b�N���lC(��a�L|I�c�n�M5����՗kd�Sp�����'��J�e���������f��0Y�u�8ez`BZBC	��&NW
����())#�������?�,�	$R��jnԐ�Y��?3|~X��ۘ���Ӟ}�b�;��"\`I�ǚ�H��(�kL�g����m8�ҒG(>�y�R�ǗIA;�/:v
�oV�Xb[��S8��M�ꗄ�i{���� ���dw7��JH$�:��Jֆ(�z�ЮPC]A
V������~����(�M�忁�Gz@�=���q�˥.r�Dk����XP�&��'���p�W5�<fl«}�ã&��������Hg���Z/HBк0в��;��Ɗ��)>]L_����Ym=N;�Y!�h>"]�̚��w�9$c�?��P�E���>`K��Yl��ou��:�H͓�ֽ
���æ��&Ay�$S� ���n-că?R�]/D�x"��d�-��wt�	&���R�E#[������= ��nƖ�[�sK_����������b�<Lq�:�t��i�����L��K+S5�o-_���N�X����P�'�Q�9���j����k���� ��	�5t;�a�ɴL�`��$������}Qի++�<��ba3��T����t�!�����2�B�-dG�y�2�����N���X�~���+c��v�=CA,L��[��'6Wv���h$� @#7�iG�:b�N#(С��zA�Ǒ�4eVB�����C%)))�p�NN!�` ��e�6���[���l�j�ު�4~PRҕ7`�z$���u{�����f� h�.[��Ha�����=�����wzr�4A��]��j�
'�M���^媘J��Y�yǻ/w�@��ybF٠�;9��^]���/�@~�*{�9I[,X:���C�&�
%���Kjd�����	�:I�%�����:�'tZ%_�$ƃKƙ	��7�-*2�D.+�3-#��l��K7՛2�]_��).���[������ ��ldX��#5.����b�Fhe�PcM~G[�&j4�~vc��h�!�P���$C
���E��~]�,�!��+\���x�9��� \����m�S�-!��	n���tP{�'��W�g:��/�~�lտȢ�џ>�����:r3��A�U��k$�N+]&L����a�{R'W�kzx�/�ί�5ľ������Q¯���5qʫn�w�V�|�H��1K�_��|s�:��Y���Ռ­r��
��Ub�\A3!�����mt�^�V�����
��ca-ٍ��A~i��L�}�[�_MlnK�{+�M$�G x���d��Ӄ�q��^}9TV��D��:���4�;˫ �/�B�԰���@��=��Ma�D[�<-k޾�>Wzm���h3<oZ|�P� Þ��G�:��#d����v��6k깾��i�7{G�-���(���A����$�$�����-�^�{O<�-��I�l� ѪeZQ _.��<8�O���Sq�[��y��{��xd��m���Uҩ��pp��GTcg� e�0��M�<v�ώ���_����o�����M���/��T����m�ڷ�R���W�/?���|!�_�(��d�;9x|���\�<Pd�&s7C�-��H�#}�J�k�[�6��!�=R7c�\��P���4����E+,e�aA��M�V
�)%�?(�_�j��\z٘0���ȰZ4G,�=W.�#��z�K�X?���Q!z��~?@֒y�D���@ˆ�+��2��673�PV9�C��ـ��t?^hw�@r����/2l/�/���t4�V��^/��Ѓu�ǹ&P����x'��9%c1�����t��3�Sϱ�!H��(]c�#���qeR�g�<��Y}�fQ��(Z5ΩOP*$��`}��S�D\��΄y�)oK��8n��ɗx�U���zP�\,Sk�Q�Bh�K�#@���m�hLr���Ō����m�*���K�U���vN�ϟP����nï	�z�nzS�o}�ӯe�q-⺼X���k䓁����ߔl&�f��c/�J8֚�9l�iL��.F|� �� ;��)Ϲ�ҢT���K����ǳs$��B-y��j�`�W�K���g��ֲ������	 yb������D灡2�8�v�+�~h�O�u��2xx�\n��W�� ���2n�!da�r5�:+�l[dH6G�lW��1Px� W��AJ����u�~�J�Ǆ��\u���t%N�U����)��U,�/ lZ�'���*P��e�uҵ~˻����i	a�=��:�Z�z�
��&}��bt���\L��B1}Piѫ,Nl
TC�)�r���b���|s*a�E
^�n�����٩]-�0!�
�ަ�+ ��i�J��c��������"o�-+�}�p�����׳��nΟ��* ��p��"Ck;��5�6ĴJt�P2y�B;o)��)�֋����@�k#����*� b�G�؈���`�N8Y��u��lJ_�&D���J�V ����÷�T���B�_ߴO�%`8����Ǟ�	���}��JR��]g���U���.'��ae�]����wv��Hp�j��-�����T$a&�o�����/��p��J�@tmb^y1n���('�Z┞�Ft�^�[
Iׇ0)o��l���י��tФJ�����s���1��9�~�}bD���>��O��y_��kX7J����x�@LΛN!�|悦��$�]cH�[%�Y�{ڀ�)tEH��������W"��(#�<\ΏQ+l&ts�{��AZn?K���<�y��p�t-=�ҿ{��L��?�b"N|8��o蟽+�'���,v&;��:�1=��a��j�v�_R@\'�?�R�����IdX��/4�Q^���/�n����M+�'�����ڳ�����.��8�8�갆������h��M�E�רyK@�$�ލ�.]��O;�J�'���&�H��KS(#\��ua3����pީ��R@)S�+�𓆉���;�/�������N.���2��ꘅ�a�1��A�ܳ���s<� �ƎPX�T������a�&ǽ7�!�c�]cr�%�e����Ǿ��n�V�����e����\v�Y�2�4,h�C[,�[<�<����^&��%ed�p��b)�c�ۿ���$�M��g�!}w9��y����"�I�簼�����'������0�������F��$@p��Q������s2�9���lK�q&�~ډ�|_gz"+������Fr}f($#�/6��d�u���%=�2~s��@ZZt=��.��0��{l�,��
(&����v��K��������-?^��7T��MK ��"	��VퟦZ�'Bv��ݬ��j���f��OIlYӣt�F�J��^�P0�^�.9wY}�b �D��_�];��&��D�~�cX:LXa+���L��a�H����NL�6����R|�i��.�Q1� H,Z��A��im�ҀQ@�+e����5�Ak�0:	e�{��(�Z!��T�;f�D�1�����J:`L�+v"]//���G�#�����'V�۵3
�p� �Rw���ղY{TC@Mm9ӪO���ݸ���;`6&
ނ*I�	(\P�g����p�� ���_�36�r��|���B�{m���v�$k�ts�����m�"������5��3�T�5f#.�.����h ���}�,A��m�L|&Ͼ��m�#�E�ߍI/^Z F�^p|�������*PC�I@�ȫI�?���ċD�1����;!5
/h�L螭��v=������H� @&�~�.�*�v�yJ�{z���&& ��!�*!ٝ<0�+]�3�R8o�XЁ�g��b� [/���)qvs��|X#3�3' �>q	��M����$e�7O˛�f~�z�Kƍ��M^¥�`�:��, ��"��9�/�c�!�K��z�ؾ�.:~*��¯��'e�]@Фg����`�r��X-�r�:y����/n+1���#����W'����'���FF牢�]!�>�������%��Oų�`b�1�g�,l8��bC���=�g�O� �Ն�=�[��/����83��'�Y;�]��	�?� P����Z_w��D��(0���aN��hGv��VG���	!�Xpd	���B������M�eB&�Dߜק�	T��imb��l���:7$���k�<I�tA��+W43(�冎��1���V�o紸�v��) �h~o��Qǝ#)�jpT�z�<!R�f�w|���������hh�_��׀�&�����`#�t�z(KIA���O��G�7�3��;����)����8��*=w���kmT�FFG>�����{���J��ې�����qʣzp������� Y�q���y�_�[�y�ٱi��vKRt�9(�G�A����ݗL�ðU�H0�w�-N���Y�T�R�ϕ�^f��`س��0��VD����-���f��@P����d����*o���6��$@'��PH��3�#����/Y��q�j�#a�J]Tь����݇=Y��k���R|kJ�I� J�)����G&��T\V�j�1��*�Y��1C싟ՙKh �� ��3�s��h:�+��R-O�v�B���K�ϡ��b�py��h��<99�����}|��-���sΎƖ:�Q����w=C�{8Y�[�=��ۯ����P檱�g��wU+�/�MS��Xo�a;e,`^A�>~�,�2��7e{6Ѳ��E � $�SJ��k|��
d�
���7���py��[�*�g�x ���H�)�~"ل��gd�����h0� �쏽��V��O�`�7��C-�M��rʘ��N��P�	�~�u{�V�.&��N_C���.��2�ٜm��Q����"�j�1u��a�P�>����%=��ߟ-�.�)�
k�N���e<��/ϛoq�ԩ
Y/onv����܎\�$��5��M��]	qq�"���)�!c��qJ�q�߳I��PĠ�s5Hd��M��V^�i[��՗�# 2�Q$	�� =@��P/̯���&��di"� �ʁ����!�wCm��-k�N����oe59yo=�����m���Udd�_�R������@ɨ;�Ku{��ve� �Ɠ��'k'E�O�J��Y́�h��U��s5�מ�5�b*_zs�<H���ͼW��������g�=��q��B]`�c�K��eF��~`���nO'i���MD�w�񃈈�t���t�P�
��<a�UCL�uq}������$6Xʟ�ے����Bm���p�︺�Ҍ��=�R�t^�5i��ԉ���VD@�7����Oa�/�PTp�3A�/���Z�z��:|8�"'y�_�$�*PA��<��x�����Cl���r87����y�;�B�(���7��;#���y!�����L��gq�-Q�i����0&B���a|��t᯾�ߏ'Y�f�vE.��`O�O�A���CmL�7>�+?*&w�%��H��h�2�(}�,�L�.=a[:�Z�ٳm���|lKY^G����
��,r%}偁����*.y��-�V�}mD%��Wg�x{��#�`�$��xS��<��ͮj\�b�U�z�S�犛A���s�$�����!���wد|�@�U�FF���aʷϳ3�Y:�,����U&�x�s$�����|Wk�4��<�|�<���9Xa�j�[12�'!��f��DiK(CsZ8c�P:��y�T}��<��qJlyͪс�x����p� �����u��ܡ�4��ܼ�-�wC*�n�����K=+��α���	��Ը�����~b������U_3���G��:q�p&��yq�u�^xj�j�	�� 4��t��k<����J���u��l���˗�d�1�X���:���-�hgC������U󝒒�=�����y8*�r�޿&��࢏��*+�ɞ�fi&f��Z՚6�X�w��Pv��i�<�}����3�� �HL�g���1avO#��T:D����S���j�z��'���N�v���y��y��4�i�wɽ���:w��W��jx�a��8�-S^ib螎��ꉟ])����]:��t�q�h=�3s�J�&�_uIY�l"����J%���y謭�����x�፬�T�����]�\]�nq��z�K�6�UaΈ��KH��"te�}N�m����M�hi"�W&YbUz�U�k��yQ�p���͋#{�'��$�����Z�/�a�,���a�C1~��	�6t��Đlll�	����%M"q#����B�X-��:�ID�z������]o�;����ş����ez� ��D
���h��gZ�SWR�R���v��gV�|����6?>��Fߓ� �;�H�>�9=
Ɯ8�:� 	�J��s����դJn2���{Ϛ{���,s5�R⢟S�?��l3�x���H�3����s���V�1h�^Ps|�ǌ\�u)�ʖ@�DG�������TW�:wG�.ա�����#����k�GZ�M��_�$�e�r]~���d	 �!��f#ΰ����pj":*JSie�OG��1�QǨ����Yb-�������߈�hR��j."���Q�����ig
b���7)�͛A�`u�_6v
�w�f�Ϲ{z�Og�b:r�fn����XU�Jc�嶵m?�KYQQ� ���;�4��,��j����غ�;�����;�B�_�LJ=���Q�̈+1ʓc��LR:�.����X:��shh�)������9�m"iڨn���?��Qs2C��/4�!��˻q<�iı���h�+īHcT@�su1�hmb�'��s�Q���Cve� ��l����v �'�t%]}���=g�.�`׽�p Ժ��m���z#˨�F�M噕v��u�Ҙ^UGeɤ;�9E^�T�%�̑�O�����5�B�<_�����9�����7a��ݨ�[������(��Hq�����.�f�4-�"�<�-��&m<��O�%�Ų��grn!Y}5T쓜|��GU�%X2�lmzK���Ne��'ÞU|t���}�==���i�G���Zړu�r3x���F�zL���MIf��`��P��O2�4PC/]�5b�E�x��LӜt����ܽ[xOik�x!��̿�cw�z�j���Җ6���P?���V�;'ޜ�l4���ek%��&W��>d[b�W4z�m�}��ow5���jDtT�w/����,�an��z�Ed��Z��~�?��%4�|n��J��	
�--�����G�w�c���K2
YIVzI�����+�=3�{��약?�"�������C2�����w]��է���x�����9+����k�?`�p3ɝ��Y��힣�c�˒����\�-��O�Zp��,�$G����Zfh�5r�����HIW�c&6
K���������	�q��kU;�~��^���Hr����CϜ��V����m^S=rt�����=7�Ru&(���k��6Ӟ^�O3$�%��F�0�4#}�l'�����������^�]eפ.Q��8�x�ډ��$�f�
������CA��,O�ĝ-kSvI�#��GGz�z)�����TƼ^D�xnK]�8�������������"���qs39%�Ɖ��⓷���k�9 !dӖ�$�u=����<ė��b���&�6G���,|��h��TB��۵��Y��PK�o_&�/&?�5V���\��I�$�ux�W$jh��(4TU�\���^�����b�.BYZz�o�f�O�$��ö��L�aS��s�B�n?˳�{5;c��6Z���̫��6wsy��S��6M K�|�Cڶ�D��ǥy��ͣi�T�F���h��UM� <�	����Y�A0�ҳ#����N�s�|�"��C2�n
𒾿�7
��MkPi/�:�6%>qw��s��x>�~����\��e�����qIP��a�I~*��U�<L6�]����޼�(���җف_;��h1|��ʘ��$OƝ9��A0��/�S�@�`E�n.����ť�U�i����W<�º�uſ�j&3��(���,J?Z-/���}|Q�@�������'�-�~�D�zu��r��w��i2,�"��g�g^0|\�ٙ����u ��z%�y Z(�xx�J�[0�މ}�wz��O�|t�T�l^�� ��xS��*��k�5Sn�)L�AE,ն����qS2�Te��<�i���X���`�sV<�K�1�z&n�o�#�3;lꯣ��kޞ�?_���.�F�vw�.@1���?��NuP��E%%�N>���5�h�[(T=�fZL�#�,�T�÷Gn����Kť�F/����:��?����o]s��~���������9��)���_u�����\�q�|>�Eh��u\L@W���͍���m?;��W3h�{�d���dd��ߊ��q�C�M�����T��vcю��h�^su�2�����<ʥ}�Y��-^6�<�(��P�;�!���v��fVJL����j@�\q��
h}�F|���E4r�X׏Ҳ2�^h���u��oMueYs&��q6]�h�qR��;��*�R����ˣHIG�Pd��`x�9��j���Ɖ� �W��m��m*&��},�BAmF�q�i�9�3��'''YK����P��{��l|�������W�����Fͮ�6����gg���������2(F���~YZ�!5�e�D6��\�҈�� ��Xդ����;t�,���:�K���̱�����w��Ym������1��q�D.�X�Ֆ��L9GT���$�s�4sݿ´���vpj̼��u뀑Jc�a̮�o��ٹǔ;<U�a�+k
*�Q��B�#I���e�UR�a@^�f�0�Z&�9	�ZT/��?��W�lO���N'~�ǧ��lɍ�ss(@���ƛ�}�����]/4Ny�T}�x��-K�- �X2�|�X�T��·<�b�̖�?�@/��l�EC�]AD��h�#iu3TrJ۬ʉ�Cc�g)�/ڊs�G�#x����L�A�C����;=e�m�M{������%%�^���K$��.��)���UaI���CS�Z�Q�8d��C]_45E�(ζ�������bQc�>5�ݷ���J~����3�>k2�c����𘲫5�`(�_�.,�4����[6|ssި�ۻ&΂k�C�Be[u�>m�gyIl�J���[5����^
E6�(����ZE�+7Hä�v��~%��H:��ɏ�ƥ�r�-�A�o�<\\���!L˜��Z�B'l[Yu/�T��ΐ��g�E��sL�>p��^{�ǖ���~h�e����5[���N�Ԩ��s�'5zf�6�O��q�ѣ�h����W��(窉���
(��.���bej�YQs��F��CC���F~c����N�Jq�����x	�a�i���Y8��D�w��wKg?P�P�qLV�m�݃��!�,����y�+�D���z�X�g���w���hm��s��3��{�cF��7*F5�9謠����-y�(T�fiM�M9;O��q�T�q3��w����vc.��9�\2���WWڿ$�T�%[��68���$��X6*�]�$�~th������h��C��/��N��*�ͬ�h�� ���2���$!�fP˘��5@'�]�@��׻�[���k	Y���]j!!��&�W��/�j.�GR��0k�U*��y�W�4�n����7i	m)P���/)+����ZTz��]�蝫/&&���揬��j�*����5���ݻZ�%�Dc�}G�N�LWg��>�'�����q���e�)oh�Kt��h@���:6L�v���B��U`"ϖ�0�����/3�����L����#��e��~&�+wG�^�ںf���ә�0iWk�7Y!��g��)����6~�T���UP��zv�\��to�6�.��\��G��>>F��}3y��ϫ����.���O��̑�Ğ#/wI^�Kÿ�e���)\�.I���]�}"H���������'<w�T�:!c�)�wVq3��I`��N�j�_B�lE�5�7k�n��t�6�"zB\����D��?�z}%qH[���{=ܻ��S���:繄	���:�S�q|�l�BD�y-�h�z�8�h}ɥ��p"U@���A���%#�V�E��,M��sR:�,�Tf�C^$�1���7���3�������s����&�[�8xy�m׳���pA�fu�`0y+U˿s�+�PI���o�:��O|����{)���ib�xwb��%�#u�ZL���V&*2g�]��4֞����~i5�͛�)�pi�� ��20����u����sZ���tY$A�f�)*��A#ܒ��Qo���~6 R�|-���xĥ���@�m[l�����2��\�ao�ی�-!7��C2�Bۍ��׾,p�'�:K�~]��OOJ���w�~:�^�:{D8�X�(�{�ߚg�|�m�8��U"T��g�,�Ƿ�/��,V-�Iw�"Z�o�kY#''__Q��J9�/�?��k�ރ�o_�-1��q��~a×��ʢ��rP�)�VDDĹ4�gM���V_�޽O�5�l��)�%��␀#�/�a��*P߰?��C���ܗ�.3hm�����Q1`A�X�4�:[��S�lll��yN*{�����/�
?*ݤ�/s�f_߉Fmޡi6BS��l�<�!��cw�n�~����\�G�j{�Ve�T�����v�ϭ����s,���Ļ��Gn�徎A�v��U�W	��$��ڞ�����sݾ��Ǫ*���&�F����x&0�!�]�P��5z����ۖvW���VZ�Z����� c�}��1W;���/���=�'=�!�ӱ��X8��m)-.���&��	�ը�hG���πv�źz����4���Q���u��q�.��C^jM��)g�r���ڶ�y�M
_�NN����604Ɋ��0�mT��Nl|�<�Z�|���7`ɫ1z���e� :��- [~���5��	�rB>N$�<�Y/��;���\ss�=w�����,g��e@��l˞()L0�)2�s��sP\���O�#�b��8�aڈ��L��G$Ҿ�&�j�d�}�0K�4���k4����ޱ���..�P��U��ۃV_v������mM�<�-�<�B�Dj���s�'�`��|��3��s��x�.5�ܙ��V�~���O7�n�����n��/�\���IEe��II	]��l�Rx)������:��NH�fܦ����O 	@��s�ޥ�78��ٟMN[����R6�9��MqyBy�����n��=%��]nͿ�6��]���ѬM�� ��U�����B+:(��##	s/�����XP(�_NBJQ���:�\����~��he>��=^��n���-#��}�=�\4���D���O������(=]6"b�!�1�� ��𿇦�y�r�>h]ë��j�_@`����2�F�ŗ�G8��S���&enz�*�9���MN��DC�/��m��x���'��?� �����ϣ�o���<H��Cb�Wm2%�e2�{�1��c�?��qmm�ot�"������{�
����"�N�d{�1Tp��Rg(�(��?��0Ke�K�����{@��&����NՖ�*JVs˒��t*�Ǔ'��2`yo�����b�cď��;U�ܴ��y���9����9� ���J�ɷ���p�KXUO�Ad{���:pܷ�
��WK�A��T�+�GE��Gq ]�����c�����G���<�g���vt��e�E�k!���s�iׇ��� f�����u���o`l_�� �y�R7�ө�� ��haN1��چ�~�j)ܯɑt�%����YYYװvbIB�m�����<=E��b���c)�rqe�w$���vFۼ���Ů��$/S~2@���s̯�Zϸ$Ґ�z���YS�� ;�h�H�8hTa]� {E7��T3��C�S�`;{�㉟���V���E���ԗ�0$�@�'Kr'k��|��l��h!+~]��'��*t��/T���>
t����%�ZJ�?"�L�nB��������h<����A��]�t�`���D��Z[��YX�Em1[z����넸B?������ݬ�9����<�;�.:�'�|<�EM�mE%ZstĚK������o^%�л�Zhܩ	��W<<�>�B�����/�I���5pᎭ���+�ާ���:�+F�y[��'⇁%���VS��|JMr�WX1��q��u ҋ���7o>�cjwi���4�wuY�38x~�|�k	�7}u�A0˲r>�fb��Q��`$���(ً�� �٩�p��<��~�(�:66��~�̿o`==��^�W9;�;�$�B�k6~zm^��˓]��m�����⍴�����@���tGB;M�?�Ɩ@!rx�)p��SzT����#o������9�" ��`_Q���F�!K�♖��3���z��-(���{�D&Ê�6����T	��oi���U�w�B��eq�{;n��!&3�
��Q��΂�w�|��о����/^(����W�z"�����j�o4{�}^���4o��g���Y}Y�V��c����c�
q��w;;��av^�}�D�����N_��豮�v�DTn�����U��m��(~
ss����{@����p�u�SKK|�Ws(�
u	g��ã�f���j�x<J�=�yd,�1##� �#.Ȫ�87�X~~~x�vbb"'���U�Av��:���=��z��ztMS4r�ʑ�L�v������O��_dV� z��Su�C����M}����}���p�/�22�P���߽{�>�x߽i�Ǐ��]�\a�{%iE;;;�N��;���=��M�|)J��z_��@���st^�YA#�Q~ݯ׼��wJO�td�-6Y�]������x�"���)c.����Dz��{W�g��Z>���xF$�aYkx����ɉ�~�PT���lF�p�G��ȁqd�Q�e������A�#�yGF�j6,I�����Xp������<>j��~0|{9W�j&č;_�=ؒ��k��Γ&��2@�OvՂ8�"�4�yw�}So?�'4�����z����a��Z�5�޻)Z��?�$�E+�g���Sjvs��A�cu_x��%Oy�������c�Eh]9У����]��;���ݚSQ�U�2�;n�3.����KH&{���Rѵz%\�,<x�!�z��Z��񩎾����u� ��WM�k�^ǘ�qȂΟW��8ha:Z::"[��k2Y��DQ����gNu_ٞ^�1>^�{�O3���cI��Wa:�~v[���ӧ�h���E��޷�O4�&������?V�dNl�-/?�����h	t�Q^>n�v��T�����Mj���ˆ��ox%�]N�mi�Rw��!ҡP<w���h������Ē�e����DK]ߢj����ӯw���n�����o/�s��ӎ�'��U�7�q�Goj��D��W�Hdj���k�?�D
YY�4V�Q\������O����[����):Z�5���<���&	����i�S�0ӻ4xk����I�M_ߘ��
+E<��g?�]di�Iב.�y�bܶ�dd����;e��;Q��c��M?����p���7o�h�NE���Nlߝ.LZ
`c�[��������F���m�m�츅X��2:V���&_�r��K7f���7r�\��(�|k�x.\UyK����˗����9䵭i��_2�ݻ�+���)n$'�,��hY�=��l9O,��5։H6��7a�F!!u�+���Tr���6�70ǆ����d�MQ �������nl�����oJz����=��_/�[[X����/s�����^����1JC�;N6D� ��J�`R��UWm��tї����M���d60O�Y��������㢑�.��8�>'�>�h���>T�3yO.<���
�}�89G[���n����P���M��1����K@�oW��Ҿg^�>EnPo����U�|b�C	^T6d�Āj������!k�/�Q�������$]�FZn���8���b��!�}}č�e�Eպ7E\��VΏ/�K�L��}�K�w��0b��l9�k��~U���rib,<9ِ�j'J�9beh�ҕ�T9!;ކĺDG�Z�Ba���2����yxx ��dd�f�ݹ�����k'd
4��P��<;]Վ"��$�g���:�g�+���öhDƴ�p�Y���b5��H��	.I���0��M���J�n�F��Z3��3M���׹�	B���&�8tX�?߁@���5r�n8b����P��v�2^HH�E��ЬP�Bi)�7�W=�;;;��Y)��Ѽ�0�xcl���ԧ�p�Y8��k��iʖ����ގ	�ro$���E���XXX�zHo���}��	pdbrq�M�+4T�)[�з�.`� �IdT����)��W1��Z86��5�
�����'f<���]B���������tb��[��*]�����I?~,,+�?����x�ݽ_�>wq��EI-�.`w9��e���;�uO�ߠ�(n[�E���r�ǋ��'�����o���=���l柕��]k8뇋���Pl�"#�!����̺m������Ĥ��w�����ý�A�[�=�m>�W]R�޶�"�.�?�����޺̹��^5X��x!V�N��Ӎ0����K���x`�v���o[\dF�x�#�;�jM�����e����jɇn���Baa{/)�b�`�:ƭ�J���o�� DJ��P������˖3�{�9C���L�BC���?}�[��廹��:[�{��΋%�Ț��M	>@e�K�T3�p0�c��}ً�G!W���ص��U��̗����<_����$mĈRٳs�o�KM��bXv!��.L*���оF�5�GXV�m9�y��������A�=n���l�B��]�����iy<�,,,��R�?6����U���zF�`���� ܫ1���f�7�e>��E��olD��T�F�RT|� �]�޳�C[�̽/�{���4�Wcq�m��;8&p
��>`��7�c�Zɫ�?%�3rPπ�c`�����Ir{χ�����ɫ����4q�Po���3����&����v������L����T��͏�Z��<�g��rmM�n��h�� ���W�CT|�V���c�VH h�Ɨ��Kӡ��.�t 	������5�Ff��fo,%cĺ�{�q�
�ߢ棻�mn�7U�?i���od?�� ù�$]�=?ݻPO���=�9�{7�D|,�:Z�#Z��ǉFʊ��]]�P�]Õ~$mZ�	��1n�V
X��K��v�E��U�4�wWF"g���~E�0�fe,z���������s�ԦvY廅��T�Gt��s��a�n��,l��il�� lbbb��]���'�����f�:Sw�⵻��k�Z���K��g����������3J���j'��8�����m��9B�@S����5�~�r�W:�)�RRR҇�zn)괫2rm�frr�}iT�<�_\RC`�ؔ�x�珻���\�aVgZ�ٹQ&!$�)��a�3�T+�i�E���Ϯ@�?XcB\%�p���=�}����i�����8�>��pm��>��y����3SıN�Mz�M7�8���bBl�����bAj?���|���{��t��ӧ��P���xHן��D�K�Pퟶ� ��@C�ާz|Bn�c&Nʮ�˸nO�ӗ�&I�Z3g�À �\}F�I�I���3RF�ޥ�x�E��3h933�u��q�%8�F�ɓ�]�)^����p�l���;��ʱ��ߤ�mzh��keꕬR�!w�J�x�#c��ϗu�?MO�O��aCy�f��a�">-,��4����卵�5�A_��P�R���5��R/��Rw{W��1��4�u	��ѿɸ�p�kD�2�0�2�_ej��䦾��"b���ח8WT�;Cy�L�ѻV#$Sr[��CK5��=�V�Y�eU��ʲl�?�h�n>�).GX�W_�U4{r������k7�쪆cȏ��ț��a!nTֱ|�����]&?_{��UPХ��~��(9�(�4���G�����|��h	�Q�������\\^PG۟/S �{ь�������wv�"M��28H���A���1{��w�!�J�k)�����[6���jf�z�B�.��\��c�Gr��ٷ���Q������ٙ��34��[��2_!�v��m}5�Q�?�?V$AFSRR�&1$+�v�Z�}�(-�EH��{��M�MP
Z��t-,(.�e�0'ot�tu�p˹{B���ݻ�Q�Pm`:""��޼�=ewU�<�*�<�ڰMNa�˸���4:2<�@��i���[-�͙�ڟ�}���$�M�Ԗ�ss�W���[�	
������Mue���s�>���c	X2?o}���@�i|`�t�=[�uv� �R�ҺF���^h��p`�7�HӪq#��r����Dc�QH�A�P_��V@�Jq#�к&�������G��);�����4:�HI�(�?*��jy��S����}�{YL>H~��i��qr�ϯ{�FR|�����hX%Ԏ���ߪ��n������8&mmm�������}}Ʈ�I�Ҽh�.�����o�`����zG�6���˗��&�F]1�v���#�W�-����ˮ�MG�c�$&O�mv�H�߫��S�����OSDzo�]�@F�'Ĥ�*ṂC�۝���Lfg�% �bW���dj�dg_���=�U�܎��Ғ�($ez?[ndBIBTt]d��6�cm-^z�Ń@i�p����Q==��w�&��TE\4�b�>wU~�ĥ>�޶�/�,����)�CF���jx'�� ����-�����і)4�_>���˰Ѳgw1*�S��J���R���N[�|����"�Cc��|Ϯ�F'[��\MB���������R��ɚ���ݗ�_��H.�=k�Z�-1��������O��b���%�%L�]��ƷKNBi�T\�S=�k�W����Y�b����r�����|%�0�UhqΔ�<�9X7���=�� �����N��v��ԙ�%k'��#+�)	@�L�ܔ�14�2��Hr��?�dߗ�GN�y�����r/�Z�J靃��k��r����%�MED�
f�7]����%���+���rG7Vi�<w(.ㇴ9��ˆH�X:;�#�{��X������#�� /A�u-��yl� ����H`A�y<�v)���v���c���1nP~���M^j͓�o���4���='g�Bur���4��4�^p������D�Gj �̒T��2}!�� "�a:����O*��/_�,����KP���Sz�'��"J�_jkmmmY�sW������7I�p&�l�$H�wU����\��ʛ�R����WGZV�-yÑ�	�O9�Y��EO5��`�8�j��KH�3;���*\�Q��ܶ�q���!`��ȩ"/�T���8�cSS���� #�.a�d�n�,/��oceZ]���F�4/��n���������O�5(:$Sv���a}��nA�B�C�a�I{^j�� �r��	������I���N�I�9��������o&8f�~������9u���U8�P��X4��D�[�6.?�J�����Y�t��2i�@��`����&ȩ�����5\�w�� S����;5T�VBqp����"C����M(;87T�#�T廉�&l�����g��R�l�gTWW�X&@MtN](�������
��T�߇���t� #9����{�7�l�a���#�B��]£����Q~������!PH��Y����k��'�=|��JI�i�y>��p��죽h(�`e���Mj��E�/0�%|��t=?���`T�U$�vb4]a:, j�~
%��4��t��#�圾��+�AR �-�S�mf�$&&�ſ!�G����Q)����]:%�VxY�Q�1�9�C�v�H�	���=���lKs��O߿ʇȉuF�߃��}��&�yi�H��@�#�%�b�+��פ�IdHSRR�M��W�Ww����W�������$�c������{|���2(R[;�U��J M�_�5L����	
Ȃ��k���Ϟ��>_�4��-(��7
�9�-����ʿ�<��M���rv�ͽ�I�
��^���`¹���n*}
,E8���)������8N�F:V�˸2
��l	���k�S5��������	�C���y��v�y��԰�GH���ɀ�ɨ�����}�^Ia"�3C��#u0��s�*b;��08����	�zW3/�=����R�ڭ���B�F��0��{�Y�|������-�`��$�*,���d�LJY��͐�����>��*K�1�74��K�|ގ���S)РE���)���z�",�~Q;��x��
bE܆��1ׇs�������˴V4b�w'�'R�(�C߬�s{��I��B�w�O�$'���W/�r���5w��y�h�k�%�f�{.���Gч!g\�C��c��M��F@�_��]e^ff��������|-B������������JH[&��u~ǍSL,�Ap�U g�vnq�@#����+��Ӗ���П������uU�cD���?\;Q G�\a�W�[��ߗ9���O��	h.v���۾�/CXE�?��B�,���T$���~تF�6��Gԝ,��4h�X��kY����D�h�M��=��\�΂�������њ4�P����	E����&��죆�u�h�n���Y����V�8a���z%� KG,y���6�����q=/?������������\Q<Pݞ��B0����I>:����#��fT�����Y'$\KE1֧��Fh��G�5P��OnUy�ڤ%-�9��Ɋ��4�=!����DO+#�0��j�a��	,�]�)�O�D�J�~t�-���`�����M�	�z���u���W�W���F �=b����D�$b���d��(?K[�0�i�nΰU;Om+�:�����RO������y�/Bc&RqL��T��^�8�iwi.�����+$�[;� 8��Ξ{n�h��m!mo޾�k��q+fko��J�Q���<;V�h	j�E���1/O�C9�q '��=ʻ=.ٸn&�������>X��r@U��+�|�9���1�vuw��4T6�͛7����JP	
�Rz����$����}����=���hR2�R����?9.��|��X�l��l��r�TI���Lb�������~���1[~ �@g���Ҫ��3�?�������)'�z�G�*ǋW��D�� @��%*���C�����^���w�����.���|ƙBA{hik�s�)~[s��3n�c���H�&�;�i�
����x�)J��p���/E	ra�}���
4(�Z��]��N�����d�r���yi�,�9��?y ���W2W�/��hDM	H�;�'��	�4
R��JQ4�ƝLH�{
(���D
�,��,칱��U���H�ﶼ�FG���ᕙ�_���yA�Z���n2��Jv?���F�z��˓�� 5��E��+t�A邛(%\��˙�i�`�L<��������A&M�h��B��z{{�hp+ّ������1��㲫��VA$�e��oC�ȈH()�?����^�	`�=�i��w5K��Raݎ������Q+��2�G��%)^6H�� ���2-\⎎�}\���#����M���z�l��ѫh�
�?U�D��+8؈�w��d�Q|� �s��"	�68ynKmz�N�4J�;[qY�]e�.Sn�aY�x�`D��*����MҶ��H��mg.�:N��B�ļ«e�O���>R�e1���:�0���O���)���
���5����Y�L�в������;���H7/�;4�Z��A#��d���)�e�8�[�����$��A)��5�3d�pps�bJ�P(�n����|��򧭃�$�Cn3���TY)(�����"�w?��{إ3�o�7Av��h]�M�������rb^2y?n�G:)ٜ�&��j
HP��}_�� |NG���X��Fm�ڧ��M��M�`ԃ���";U�K���ʪӧw#l]AOOo�hgJ�ځ4�����L_�>1ؔ��]���;;\�D�X��ؓ[�v�h�$����.�1��<s4�Hj���>:��3����Zp��t�2n >64Q9�j�ϵ껇E��\���@� Pf�A*�} kxm�mH��m)��$|]]U�>�N�\	ݦo�Ő�'�~K�-$ `�fͩ�>�RQ�g��g9��w�g�`f
���U@����D�Q+++�M���%�Q�ժ�h�h�p$����[� �n�����G<=F.0WGO�^��ۓL�u�߹P����i�l?�#�=���	��{��>��Jk8����M�D�x���}�up�1x��Y�xA�s�$s�f���x��&�W,������E�>��>V���[��h@��ᡐG}$��kE��}w�>3�Rࡑ�M�t`��eL�$�!�&L����wZ���7���L��d�7J2��7b����N�+������T��2�*(���e_B;�9��Y�H?㜦@�𚛛G��H�J�����CiR�3K겝�ү����fgAZ��ZO�I
�OK���[P6�&(A�b]C���yu_غF��tL}�ҟ`�2l����W������`��rGQ߇aB#������֍:!j��w�beܑO2�3>iQ����7�4%Ѻ��M8�︝�W_0�2ɜX�G%{�F/�a�ـ]� 8�Q�����ӓ>�2����kA��}����6ͥwf�J�f�����^�\�>`�����+z߬nD"d�>��N���Q
��.�z�ѵN����a�ԙ��[�A�X��Vx�N�d>(q�j>��+�س �JQ�4d�J�"M�~�����~|��8���}��Kc���A@M�n�ؾ|y�?���Y��~R�)�<�R��s�9�ƻ	��Z�I;h���Jϔ��&^�(U�L��O|��&�ϯ��/�ۋ۾�
>$t�ӧ4��E�­b���Z-�y��
����M�+�8pS2S�����V�����6�� �
�	q�B'����3�cX%@��F���u���F�ZS��JƔ]��F��l?§�r���H����Y^���O��cN�sg�"l�uh��]m۬��"C��8PAq1�e"����6�M�>�J0V��o�S��''��d=I��n����@��#䝪��G�pto�n��wr��l�>���F�(줞K)����e�g$�����^$ڟ)��x�9;��K/��	9%}��Bޤ��SpLN����2�\y���gf��>}z���+����ן/Pj��( \-�/���Q�5.��8�\�vw�^pJ��#�q����7ӚO�B�s�v٘���PK°���}��_���<B,���F&�C�����Lp�Y�Lv��ڋۿ�" �"�禧���@o�R�22�|"��9`���$o|HpK*�$M�v��X����$OrdK�E������\r�
DZ2�Y�88;������ ��S�+Wl�:�?�]8_��7�����C!]�ZWG�?<~��?,ɝljFw�M�����5\���z]{u�M��f�53���t����;�����Ecc�S��r�S��ɿT����w>�x=�YU~Vn{P��>�K�	5Mާ�AR��!�c�������_�g�ǝ�H��F�h�Bn$q a�W(@wr$yAZbϽA�7iiZ�,�d��į�]���������,��k��O��ߜ��w�'��d��\oA�����R�y�2��;�$�����Wf�K]]����c�#��0�p���<N\Nd����ϟ����5�.�����4%
;1)	��w(#�i=c����l���d�A�9�b7YXY�)��x�01��!��]���4��4(�#OՔ?b�?]��\q�E�#�PJq�L;� Fy��(Gh(��p�ϴ�x��H	q��[�O�7W�*����#��C	��ݣ�¤Q�G!d�U=D�eX�Fqy�`lPSQ�����r9ƾ��9J�ƀ�xǤ���n1i���	-����;s�W�:�G���9	R���^�s(��a�k�7t%k�~�Է�X��(�t�J������r�����)i,�gc.��W�9N�dwr{R;�>>�u�))�@<]�F�O����*���8OqIɝRО���n���冢 d�Ǧ��䔐�pP*Аb�������N���@�����}�%��kkkg��NGm�窭o+KK��RT|�]PP�q�LW�?E&Se@��2N�9@!�Meʭ8@4��q��z�e�����ى�}�v��>gB4$��+-����/��j=����������f��v�}qĚ/M�E�������<o�e+^j�͗r�ϟ=N��������?�
�������M� G�U�&��
�
9��Mj��>���}-s	�uM[\��XE旁�����n(�V�)��N�W(�ފ���f�9͉̈́���'�|:�t,/ =p�	Ў?Þ�:+ū^�q�h3��>2�J��VW���X{{�l�B6��CЮ�7��]EjmpA��Ii&��s��bTgڟ�Ƽ��������?�����.�>\J�}x.!��I�۷���i�>G�6����x-Sz�>�H]߉��ݥ~.���KCa��� &&1M[�z%��9��=�bbu�C9���o0�>��$r��75!_�l�u�I2,����rN�������.�6{^$�*3�������[Ʉ���j7��\\�q����͍`yLg��T���~�%RR՛���L�wA{��z���ϱKuw��MF��%���n�t�(�Ң�5�0~�B�� ��	���PWg��Y�U���@�s0&�܀@���"Op�"�c���U�����v��:���&��� �`H/��^�����h1��'n�@>u�?#EG85�g��	ص��|�'�g�s�gh�(�p���f��� �L�%���t,7uS�\���]�%qPB��ٳ������h�&U����,G2�
=��=/5�_�o�l~��P��@�]mO�#�>��������Dj��[#� 1�i��m'''-������D9��N���7
�$�K��׼�����$	���ԟ��Vj��
�j� R�n�UvP_}=B&�1[�S��8h���SO�z<D��G�~��HIK�* ��=J�L�0�$�Aٝ�YR`�G
�Ke�70�����#�8*8<���}���* �4� �����a�=�_3�]�9`>ǭq�h�K�舺��K�u���{�$y \���A�w�Lq��9
���_z�&*�J���4bf8C�`��F�[H�S�-(I�D�hn��P��(=B���{�<mW�����_���=��WT\iۙv�MTeK��P�7yȫ��Kם3h4�o�o'�kN����T,���.��Cϋ���Mn;�r�p�o F!q\||#�e��Em�\��ޥ�C�F����,9��>��S_sJb�?U�۴����)ߐ�j�5��W'ud�(I%�[��gg�H�����ZM�>Ai����W�m�͟�n����>�o�M��]�~�����/�s��'p��/��'����-D��ƃ���+PZQQQ�)�쾐Z�8�ׯ_τ2F�~z��>����r�eA�:X<�YK���6���3x���{u�:����-j��7�� ����bo��jh�b*B\Z̘�j-9Xr*z����hG�ׅR�&>=o|�I�t�	\W�U'���+W*�4�������23/���y:)JK;�kh2ƈr[;m:���~�3W|o,ba<`k䟆��������*J6 $)��Dv?ò�O������W�4焆���Qr臮�Z�׈��*��2�����p�1\,����Po����<A�؟��載̷�G^�>�T&yV�U9�Kك��Xx�aPƴt�����:�H��	�÷�O�WW���y�xߞ��������^!""j��L766֏1Z;!!!<{1��-_���apd��'+��[v�)ǜCŬll���t�
[���@�K����*�eQ
�>=�����n.���.��k�Q�222;�Aj��?�����\Q�W�x�~�aĺ}��9[Y�	�~S\��5��e��xxvֈy���������k�`��;�$ZE|�F*�_zz�¯��t��o�|
��!%'�'7j��͚���0kӆ#з������x�| WMMt��ә*Գ���[[!ZE2ZZZH9�hU<�������`s���Zm�%��npp�����n��Ga����
/�*�4v���g~����M�i��RaA��fE�Z���������䁟?%r7����u3
Q���!%�eIU�Z���k�U܀r�*:�(��hw.AA*ȁ,Z8ծ3��`�[ P��b��Nh��f�8DMj*wpr��j��E�j`̖�uRRvc��Н��ү饞�C�eN�8����8��tY[H��i�3�/4� U9��"e��؂�����CE(x����B���u���"���m�V"�?����#��������lF�L��!|a�=^#N*N��w�]��w���LV]�a���p��q-�f��x���d-Wt�Prς��Ǐ�2�पOv�K��
�ݽ;Ow9��|D6������ZQxcʸ⹥e��tX萯B����2S4��E	k��������=�������8h����Ϗ^x�f�T������dd��+�RR"�|��>H��𾬬�`j�1	��g����;��y���k������p}�䝋xv����-w�2�0e��w|�%��LL,��ijn�!��B���� �(�S&�CE�H��Mȼl�64�k
���vh6)��G�y�c���!�����+B������]Vde�B�=CVB��P��(�d����u���^������s�뾮�����>�?TR��\�ؚ���u{{^�z��<x��Iϟ�޽̛I�2�R��x�]c���y�vr��T�I7�Oʇ|���Tml8���&&ʼ���� 5ԑ�����%4s=��WRr�b�N��/�Q��80��-�Y&�~)��������k(�� ���1�����%��[���"Y�r�z{U=z���7D�]�u�-�mε�2�j���2�|R9�nݺe���&)+����Δ��\�@9����ۛ�Ƒ�����,P����s��>~�|R�#Ny�I�ʭ[T���XAM��Ƽ������@R�IR""f?[�d�a����J�i�u<#�{�n�E�d�"[�N���{��ҷ�#�І�pT��=�[�
:�JM�$�A �# �/�Bxa�U�G�n�`aa����	��Wf݇�%<�X.++����9*�磤���fK�}���y�*J
�flM�k�R�V������A���<
�
�!�K��L5�|:� �����yysّ>�0���R4��4.3�r�!Tk˛#�)D�o�훜$��!�4,��YTT4ͼ�FgC�tt���թ*
qc��>�V�u��!��׶�*��'Zx�#y>�~!���NN����ѐ���10��=2��̠����|��V���wj�^����vlZ}i����8	OZ-��\%���WH����E���Ϯ�����R�i*�Br�}JO�l���B��
?
�x��������1/��cN=��1U���vU��T�VuMM;D��P|����ׯ��Bxg4���CUy��jI��	�o����Z�w��)���҇�!��a�\�w�Ut�U�����RSS�	�Έ��*Trs������zKX?A\8���j����$ۋ��j��|(�Ш(|��$q(SSSQii��,���rJ����-�,&�`T�%�C9���U:C�O1hK��w�șȹ�������<V�J����%C��S�����������u�AI%$�C�������(��CM�\��"tx�4��7q_?�Z&��=[���RBh�ǥ:�	xP�<��
����Xjǈ�۰�;)�#l/�jX>����Q�ƥ�ka� ����566&R����OF~�!���[�c���od��l�^�����M^���TY�->��� �j�%R���z&&&����ꆚ:)��d:�K���V�;�WIq[���n2�8�����/�T�y��XE@[�∁�0G�п� ��q��}��Qqss��;o^AC~`�aN�`�ޞ��}���H/TҸ,3	P��|�����P(}�?�O&�-�^�ꨮ_>mE�����p�1n������;�x;!ee��wH���c�oH��45�'J1����ݪ#ի&`�}������\6JJJ-�����yqO5l�q��M��l1�B������0
1���5O�~��"3�.����.A�!P���r�/�/_f�!`қq�6���M�p�����3�
J��rCC1ќ�v�(��d
&o�MՏ�?�@���&����u���+��9���W^E����̗/_��A�~5��&^����[�в�����P:�[�SO��f�>>�[
� ���Ah�Y��/M��<^\Z
y�N�Đ?x��&��Ǐ��:7�(b3�?�ܼy30=��}��HEUu��{�����������(����j�����y*�����ѹVu�РD���
�VӃ����\WP�x�G���ߏq� -�g�A�L\�"�)�PX����TZZ
@�����JZ������m{5~������Y�\���8�3O\ƙcnݻ�]j� �&B3T/,����	}'���Ԁ��?2r�b���������H��93HƧG���� i�|�I�!����/�q����KKc���j���Q?�
V�5�j��H�V�S B|�b��� ��|�S8n$y�@���K���塞@�`��u���QG�?w�--��K�7Wi����"������UUC����=MI	���E���%����e?��E��{zsj���5�+�&R�w.��<�����Ͽ;��' �.-���4�VP���ͦz�J.���Rrv�8���Y���w���DAIAwrf��C��g�k~>*ʎ�����"��odDrɽ�/uFMm�E�4>>�+�Sԗ�5�Z�G�t;{�H��r{�<�vMj>>�:�~�-Bb�V�-�kT�� �g���q\�,��-�Qa����D
�\��ދ���v/�����I�\'#t@�K
��U���"�GW���9�م���G��?�TA�F#c�.3�^]]u�-7(�� ���8������=�6�e�����h�v�����\��A���	g���k��Z���u޷ �>I�������}����d�L�y��+���D�b�����Aω(p�^a{�����,���`�2B"�;vv���-�ܯU�I��%��p���N��?.�"6��l�&��H�Rl???ZF�8.9��B��.`�Y��(�A������ڿyC�����Sc�H�Y����͖�W��t��,ԓ��M!��>	(+��j��zF^@͊���������;��}����"�����JI;;>~��(h�����k��t���h-3s��H�Vż(�����.K�;�f.�|����<?�����W�L�jW�4���߶��SW�b�9��&Jg3�l�WLL�/p�2{*�P1,�`r!��?�)�s���]����û����w����	$�L��`p� �M� ��|��H����X�d¶�uc�mc?<�{�E��2T��H�� �Ʒoh8	@4���D�!�V�rY$�)�#�>�y���<?[�x�<˓CGx����,-P�UOP$��z��~0�Т�JR�Ka�)|��[�q���G�3�$r%{{ZwXO��s�
&Xy6���- �s d��h�#����	���9�\ _ ���>�$�y��wCT%���h�?��~vYLY� F�%�t���?���?j˺�%ϊ%�I�q3"�z#�g�<v�k�>2��P��F�<M�(�0�ckq<����,i�+�>B6����P���,�{籱��G��\/�x̡#1��w�.k�R²]���=�2�i��/�ݻH|\���:vh����%���p��A��N�o;��|�9�g`gs���-�r�����"ސ��Q�/��~�d�B�����B������y�0���ZSc\�}M(� 2 =	���h./�3��+BKط��p��i%�N�0ؼ�� E���O��e[':���\p�j}�]��|
�ې����)	J՟���6��f��2��	�]��	I�	#o��fPb�-́ybPBt�RO|�w1X>�A�Yi������~GV�&'{��b@��piB̅�KHغ�V}x��
���k��P�{3���LbUΕ4��h�Ԙ��	Ǫ$G6��W��;��Dr�ǉA̚@��t��'�<�����w�I��3��""803d��t�32�kE���d�IqCT������qMʘ���>�%�6�⯆�_{L{4Evh����}�V0d8(�6I�_[�L��ӡ���e��pe5}�(/4^Aơ�8��lml�V��BHg8��0��(��i�(À�%R&pĪ/+E>�yDk~�ȿs�72�����d��c��{��[�K��MMd���1���m��jhH_��S	I�U9�߽s�:f�>�N�3���Vs++MU\	f�P�_�OH����윜lhQ���<�s	�I������u��h��ZpEW����5������=L�diU9�a���iL$>RFZų/& ��_R�y*)6��b����<���)��1333�T��IO��Pi��*z���NτT����\� �b�/"�4��9� ������.���w#�}@�NF�J����]\�K�)8q��u�9��֘ -��L�r����!��\�62w5����$P\p������[�ڑ�(��c� 8U.ދl=���5�U ��$���j����A~]�y2K���z��ctG�|�W^.ĵ�Ƌa_DKm�����h&ޚ���)@�^mm���9��xx8��1�Y��e)��q��x\�h
P*��TT9EE<�3�y4M!e`���^�X��X���ӗ��~��5�3�pN9V�t-�o�bw�㼤��fv����:�6?�[�A����6&3��%v�[M��ZC����sww(�L�e�V�9�鏫��X(�B
У�;�B��e�N�R?Ev���� )��ө��V��-	�����%�ٷb$X�d�����"
�7!�Fo,�^��� o����۲���a1N<�O��X������NvI	�����N�=��Ks�����H�]
��y��T�o�,˒g�������y���qkos��J���v�0���SNNNv�����8M��6����F�=@Ů�D;-�
���[?�<��`J�Z���]�yg�'���L���K���2�� ���/Y���8��R��í� ��5qLB���a����<�2d$m�����W�L�}
mV���ߪ�w'��B<hc���V��ި5r���`f��>=(�q��i�s���t�Y&]Eh��ܹJ8��I�J�&&&�圠�E�A~�w�Ҩ��<�������z/�w�Q$r(��zk������[�,�b=R�:Ypx ��x����4E�ng���# )1N:HSw��Ǭ�������A��{���ʘ��5?�7�7�M]f�H��"�1^7x��|��~�i
��!)L���
z�	/T�y:N6Н�4����~����uH�:#�~ղg���� 6w��������e���p���=�	��	��5&[���*���6�X6\u�)v(�ӻ�\]�>��ͪ\Z����	8S&>�]�CH�ݯ�fT200�+J�rY+���1+*�:\��{nh~G'��H����F�$��@�"~�����1��4I��V�a�{�v�����76T��$�Hm�)��h@M�_t��Ԃ�#N�,���� 3IW"8��hh�Gpv4e\&���3??_w0��~��Oh�kvN��ޚ��EjZڽ�p�B�G��R���..Vps�bm��D�2��Kc�廷��mbF�����~,���'Zh=H����da���C�����k^I�m��D��t�渲xJYcE'�Fn������+�4��*4���scO��!�Z�}���(�J���]�ɵ[��j]:���2^Ȓ����?���t%�Uv2G�7w��V����KH�(�|	�[B��h�E�]�h�Y�h�5z����q�D����g���C�3֝�Pl�6cb5&�������QT�o��c?R��~�{� eb�៫X2�D<d���'�,��1ui8Y�(����RB�`�&q����i��dM�v�zF��t��h�7K^���zQ^\�rץ���Ӎ��H���zz�I)�!둵��%4e�4��u�X?�r�?Y�4l���X=E(��]���O�&]�h>;u����^�`�%Bh�sq�������?��O��	isg��kɬ�SRRj\m�o�4�>���6�a��"��*���p#�����$�f�2�����N�S��d�0	�(��oL���e2���%�ߴj��H0T�Q~�X?��5���X�:�]ͽ������~���2�qr�� ���_��gh��f�2d� �\V�{�|��n���3����J��'���煽2�,+����pZ
Q�!�D���5?� }��"|��Xt��WOp�����U���B1z�4�ϬV�����og{C�7�\b>���Zq��b�Ca���J�~�6�r��u�^�"�����S3�q�[6��>��m�e��ݻ�*����Z	K�������6����/{�3��Tt�W4$��D!k��Ɋ�P��� Ey8�+ikk����Yq�exg��-��|ƦN�4�$�o�j'�{�5>M!�=�\�Y�p�bk	r��N��0��c��/(��q b�&3O�Z�TE���.�����d2.p-bx$%i$�]��ȟ�=���ܑ�p<<<����j�
�n[r?�/+�K�b~M �p��^o�|�߹���߼�b/5�Ύ�ݾp�h_��}�	����o���(�tRRfEH�F��AcNm��p뚏����-��h�^�k}<x�	8D�I�����i(�/o���=�^G�R�!��,JKX��yv���0���+�|��1�x���	����d���,ͱ�&����/���۵VX�D4��VLl����~�G�~=paE�g����uӥ�:�N�E�¯_�|�Gѥ��{_�c��6�f�����.Y�10�X���N�~�MQ �����/a��-ݒS1���/99�����F��)&?�%px|~{���=USS�gqɾ����o߾�ן�RF(��2?�@T*��#�E�f`��G����?���\��ƪ�ޮ���>Ƚ��	ﮌ�9J���p����f����l�e���pD2D�� �6��F;��0I���U����`jtIYY����k�n����W���qh�U��bEҺ��l>�,�mn����Y�Ym3-b���0gx�ڟ�߳90]o��;::�����BӴy>qj�B30t����~�q�6"����7ػ.g��_�������]E�k�$�Z�$��W�C7�VU�	!P�6* �c��Ç���=�F�v����v�Q4�}^�~�7�>�)5����G����K�ɞ�J*�8=��?��'k'�p�ݡ �=2��x$�r`>��G18���x�1Ra��ٳ��T&�&���oE �A�a��T����8�4?Eo��?_�^�!w���������KF�s-⭏?�E��-��S;���?�pZ5P��UZ\Q�����l���j��$G�V�[�1�Ai�m���ׯ_U�(N��c�]uf�v�����Mx[PO���6��o�>��O�j��������O�<6E�pb|$h	� �G%��9Փ����Cut��,�׭���<��Ťu�]q�\.�b��{�Ifv���s�g:t��=��	��>%^���&��6��,�&O�^�������\�y�9�
�ʈY0������cQ禿���∤6w�޼!mp�Vs��]P24��/�����>^�T�w�^�:�tKB �����'i,�O�|ϗ'a⃌I$�������f������z�F�{��q����{Y6'���#(<h�z�o��6�.�L���+M
�Vg;�Q����������k�ԂBe����������98���$>F�`�(l����I�	-��ᡮ�����ޢ�޳x�TתF���\[[��n�����RO��9�����\C�+�%p��Fw�JNJ-�2�4!I�������Z+����D��G;��nGk���\�WE?|7�q!��\I9�&j�d䕮k����0���]�4��xxy�T��.ކd�PJW(d���&��7=���g':)IZ���	�Y�A'�\A\A��4�i[nY��n���}��↳���Bv�z�F�F�pSW�����f���4�*��l���dl�}�"ͽ�\��������`֩�r����0;�����͒!>�ԝ��d�,������	���6��QM T��wS�~��Q���~M�q읓Y=�,I�I��\iF�ha9��A��[�bbbn`+fc�z"?$'S�y�R���@��S�:�(6�����ƃ����se���#B���7��qё\��}=�m?T<6n�y����.���R�-�f��	O�I�<Z�TF���pjL����Ĺ��Y>$V�B���N�3?C���ͪ��?�ehd䌗Z��ʦ+����&T:��D�Ê"�q�!}SS���֖�ʒ������ ݙ�á|���G�N	,���`�_v�ɒXR���� ��|6�l�.�-9�X��ѿ[�	��K���:q2x��N�K#\yRP8��������1���n������a;񩿐����qG�OW%P��p+e��n}f�G3�.-/�O��L�� �U0�4L�E����l�LM����P�x���̱į�S�R � -#�'����e͖��W���;�>�K��615ퟚ��L�E�b"FV���2cc/ӵ[�i,d��ʟ�INz�}�ul���ŗ��D�~�oH����8��2E��� ʭob�-w/����&x�/�����F;T4Rk-�o�$�t����@�u���&�jo�T��C�f͂��zۻІD��B$q��8�N	2��Y\i����VV�67]�0�Yr�VʋF�A3����r	v�����Po���'�����N666�o�(}gJNMMum�2���)�$� ��ܜ���V{K���4��^��)�R\��y���qW˲~b����8�=I�ng@���W����＝�c��';����vp��B(�,'D�[# ���*A��K�OB�8�L��5Z�I��#ږ����gq�b�������:_�m�����P��W��dd�2k�~���Zt�Y��ښm�Z�u���2���N��j��w�-�/Z��VB~3�g��	����M��SV��	�B�Ҝ�Ĳ���|	�rw��#��T1�Vsο�
Cv��-!�B��t���咊8'gÒ��a�v���[?4��P�t����ڀ`(�`��%�Ɯj�g��j}�VD80F�η��z�Ǆ��AV��>
����}}o4t�.���-6t���{�v��+(���	������Ň���N� }��!	�*N�1��u�E~y�Ɓ���ŔU�ެB�"EY֘l����DU\�t��iQ��Ph���w�i_ț	���c䶤�a����2\c�x�Å�ۊz��	B!-J$�B�H�*ώ�n����?��t)����^Q]� ,,l`�����_{qu����Q��_>��ʮ�N����~�7�Fҥ��j�,�JJ�1������d���r� s�M�j�?`j��'��7+[آ�Q��?�����kVV���#๯tl�up�k	Ė�(h�^SL5<�Ņ�����4��T�����F�o)�<S�kqc�3����������qr�v��$]:����+6��O}���ێQRj�@�3���ϥ:�M8�/�c�כ����I
'���I��SWS��.x���`�$ "''��Crxh�����.����u�xW�v��+�y:-�<�JR��&�M�[�]�v���cK=}ABBb�1�HKK�%�Y��� �;\f�D?���El,�<�PF�x���L���;Js�5�����H��?)*��i�%�|�������� (n���.�!F����ބJ���++�d��	I�ތ�C.��ޙ�������߽���	3UU4:�\��UO����p�8����I�{<�\��e9��~>�2��e1���Z:��E��Pq�q�*r�(?��hS���95I�}�������ݐ��3֘�S�O�B�{Q/a������M]oU����c�=���H|ٮ88؆Έ�^\��ۘ���#���O��~�
D�P��2�l$��/���+	X�o����J������ӡ������i�r���$�>#R���2�4�����w`O�z�z(�@z6��eݏg�Yf!��W}��gK�z�n��v:����P��DY�r�g<���6��Q���?,�j�d�o�����A�K-���bP]|X?A����A��g�uu�Ѵ�,�k2����E{J����a�~�Jy}��}��]Hצ�u�!��e��m���sr�v�~F\؄q��ݮ�%��Ƿ�2�J��r�&���z�����s�[*s�Ų�2;gg�z_��@�[FC3�������^�� ��KqNMMM�IϹ�Ď��+e�|�O��ⳎqW���=9i��3Dڥ���]t�0����E�r0��`
Pώ��L�3SR���^f}�ȊC-`ȝ�=u���~J�����b$zo�S����j�l�bW 6��A�t��nDr:%���#�R�o!�0	%�222�=S�<B���L���L1Nc~>���=�����sF#}}�Z�y�%%%��P
(�Ės$�٣�+g���Lצn2X�濚�[�(ꦟ�%F  �b�7�7�\�eȸ����i��c��(���o�:�
s�/�Bl�m��Nۚ���ݻ����W�����<{�{.6
/�c���J��I��7��/Ϋ��t���*W�\��v�*����_�'/Ǩ�A�ʞ�I�V=��b�͟�����#��w���qrbb�C�{��q�g�*��$ءS�v������D���Y��Y��&��h�o����{p�q�\M��
jԶ����ᗲғ�9���z�ǅ`���Ǔ��5k:���塒��z�Ⱥ��w/66�����m�S��	*��#fcg�;l���v�tH���aې�����{UF���f����k��T
�k<�SLȏ؃Fem$��)�[nԡ^^\��D���Ӌ�Oz��
F���C��bl���edh�\�2}�y�u��rCfw}�H�!�P�~����a4�	Uz��Zl�w���g>�$�t�)I��g�%�ߧ�y���I�Z�"�l�[R�_X���-4�[nCRBB����Neu��6;j��p���Դ4�����Ol�����{���w�(sV�![�Ѧ�, @tV�����S����~�:�x�6VJ� _cִ��(�O	���1�`|~�ؿ�`qD��'�a�@�x�{yMYI���>²V�!���,x�l��I����L���U�O����Lk�S��ˠA<���,��t2�
���G}���F�r�b�?���IYO�"]�^���:hhݽt����#n�
'GG3��g����y��^�O�o!�b�YjQ���9���~j��,OԖ����g��o�j5��A�i�r������@�Z~ˆb'������S�s��1v�?�1��m�C�0@�Ox���c�����4�.�f����#�<�LZ&G����Z2��')��r��-U#��.�;`��%��:���ed���t���䦒�����ʢ��D���VܹAd;]B��~�i�G�FkL�&D	�lہz�
tPƤ�|)��-�hkk[��������Nz%�����E*P\����ހӇ������x/)���\�-�ȑ���^9�wK\_���M�>���Ƣ!�s��
>BeY3�|U[�W�Q�������oVr`�!B�dL�Ŏ�u�<�����/�I����S��XbRŖ%���F&�J���F����{3k.Ѿ�4TTTOm�|�V��U+k���?���� *"B*��5N�Ug�).!������+�	�Ht���Vt���m�Z�A���_�p֐?��$wh&���s}[aD�G�|�j���w����[���QHD��@�V8�$X�s�M��			-_i��'��~���:��N�.~�K����_hƚ�SLmXD\R�>��mvK��' �C���2S�v���b/rs����B��Yτܛ씸fba!O�;�IpX<��Ӥ݉8������_̅����Q��
\�h4e���,�tk��$A�A��z�9�al=Wǽ�����j߇�`tH6���D�5#��@�K1�]Zg�'ȱ?�",.+��Q����^yy+?iM��Ņ�q���M�|fB��}�K���	&�"g�Q&i��Pʣ������.��Z���vww�1�<��%�5�clL�t8T�
Hrm��i��"��A��Ʀ��s��0Ɍ���"��� ��,�u�u�UhU�r�=���g�h�������}��[��!�6�K!��`}�+cbm�HQ�¦��ZHZ���OڿL^�pt]�C��ӣU��ͦ�dRF���V��I�#r��ȃz�����j�C����]EII�Z�`��D�J�����5�RM�^�~|Z�WX���Á�a{��6�C��B�9�)d�#B�~��,?�o�y�d���o�k��)l� +�azD������Fh˟P�	���_�0L�Y����%"":�R���M���X���!�oPz��h̩]����r렋ZK�p��=��9�|��+Qˁ����@c]K�dR	i�w,-Q 2`Wv��r)YC��TTU/���c|�������\��Ujs�~�S�W�VA�%�1�uI�驽�(b��G��K����B��]ɝ���	8�h�Tĝ�3�t�����h	��'z���b��u�}� 3���W0�d:��l����Gk]X�s��%@�Gܕ"�jnn�>fË蘿��1�P����J$��۷��Ґ#u��I��+�%������K�'Yg���A���ed�����x����V��D��_5�C�]]�8� ����n���`�˱��T��;�{x���GEx
����^;��R��	
�+����I���W+:5���
���Y�A�~c��a>�8CFiO�j�4f�d�/���^���h����6�Jd�Dy��� ��ތ�!{=����b���H���&�����:���IH*	�Q�wtt���Y<@n�,B��h�����<}`rd��oG��(!�J�����^�%TY���5�ǯ�����6Vŀ@�sOϩ��P��������Be0fz�!�S��ӗ���_>-|�/��f�.h�.&cr��L����Φ�t�������2������>�Lh]�E@�2^��#(�θ��?������i�͏�mPo<V�#p�_N�EE��&c�y#=r�7�ߍ�N���7���T��m�S**H�+$'gn��f�k9�������l�����'�(jĶ��IY�eQ�\/l]�n�츛��wE�O9V�<Aj���,Lj��r �p6L�:+��n�D�y_�H�������k���˽���鉚�<�����6�uPSR��@)�Z��L�#�+d��ϸ,a�^�w��V�=9u�2%��Ѡ�����p� �"�zvMT�������r!/�',���qdA��O|�j�o�t�ױ��5H�(6B̏�������JP����(1B*�8
^R�D�0\�jy��Y���ٺ�����r��L�k��T�
j�������W.���1ה?C�2����GSF���\V���x,|p_�x�جT+��O}�����3����`��F8���1�R��;�����w���-ʋ{"da����jdaG�8�m�d��Pgf2s-د"�***�߲(�s@A�O80!M�Z<�����y��T�5
�#�����x�pM�9�F��~�+����$���4�s͙}?b�7�Z!�~������*Z]� �gD��L��?��w��sc2l��(*�gC�А��<!�S�h�1�Z�X-+�V���������޾�#6����9J�XF��s;�½��%�\�gE�q�~�m�X�?��F�*����>�&�<��Êl�s�h�_��ŃM�����ܹs�U�H@.�Ԙ�oJ�xYWN+%�e��d/B+�=C8�*��MoW�����@�����%l,T������'9�j�͇Ŏ��M��	�"��b{z�Wgd�� Tx՟���h��Z�-��f.u����+����X�}��lqeEIE��H	����^=G���+�M���h�����t���h�����I�`~KF�>9���k���'w/���lS]]��֯q[5��{�*m��ý��W)v�e�T(ǎ7��W|���x�7��\�#�Ǘ�}W+#��z�	�څ_�+�{�#�#SS�w��w��E�~�Ix[���� �|���h;��g�m3P�{F��He\��ٙ�d�\g�����l�`��ן��o,/C��=n:4�@GZ#`�:T�T��l#����( ����"5�Ϸ6�1����MU�2�[�����t^��Q��З\G�x���ם������5M͹�׮|����/il��e�������GYYmjj:6ږ3Q����〺��~,�B qrr��R���2�l|�v�X�!��j�q뽶�N��t{��Fs�/C�;]�����(Q^?n^�g+nt�SűܫZ�DD�-�����ɖ��Fo������o��fͻ�*
���vU��&�_J3�y��(�������Oc��*�py��Yp�}Ĩ�y����CII�����m�Q�F�gW���%p,����tV���{p�Eٱ���:�ݏu�ۇ�)�?���!췤.��Z�mU�m�B�] gI�����_ ���圇���g�iD6*~�����Q�ϕ?0=G!�Tϟ?��8�lPfr�d(
Y�
�1l��p�NI.X��z�=�80
n�42�sO	P��5��]���_VZ��XC�R���3��?x�&��.ks�ܣ�4M٣���R	K�&e%_��D
ԖZ'��I�*'���fff��\U��<!�0P((d�mp�B��;G�ӽ��N�S��dSd�{��е\g#�{��o�����o�ϭb>T��v��B�H����J�E�DL���"�'4�����j�ff�U�	����VGg'�4�N��+A�ݜ��#;��֪j�ԋZ�ۭ���j�fgF,n��e� ��V�G�R�{���^jYj�����1�f.5>�{{��rz����&l��t_��I󖎎:����7��m&��ϱ/R`B>~�XTeʫ�˱؟�@ixmUom���ϔj/*+[:�-,,���	I[tp�Ґ:���LS�׷����y�+
$d�!���q�� =B��ҟF�R��2N�y�^��e��6�������;�NƇ1��_��z.��ɬ���a�ht0���.�!�h��v*=(L�[�����**�ʸ���r{3�F����+d-�pO��xv`����\�
�a������'X�{�DG��*�ٿ���DnV����|�=�&��6�HE��[.�d���m�[V���V�<��F	v��W�.��L�R6 �"Pm���7�r��+�+���n/��G�����W֊�̖���Wܼ�;��f�{�,O*Y�մM�<�V�/�\aS��3V�5�Z�����Շ.��W�>���}q�����>���X⭙�#ڐ��'C�C'����~%^==���z��]�g>��o�	����D��Efo�;qmt42<�Ns��.
��	��(:����(�|��O�<���k�Q��z���<V�^L��W��׎2_`5~��HC��̟	���T8��M\�,t��*�_H�o�������^��G\=��ꬩU''A����Yt�Fv�A4��Swjnݺu ���{_�\LSk�k d��]q�g�L�B��(udZf���<M<�z�W��[MIV�]ɂ�F��XEX<rw��V'�Sz��o�hH�(���8c���.=п�����I�7_z��bq�l�|��$2^�l2���x�ki�=ǧ�.	D?�zyz��>�}�"��ģ�6[�m�U�R>>5��Zk�4����:htH8�kzL�c��H�m���K��÷}8�< �t����F]�z�so�����`V��ɇY>�|�6
mY�%Q��hᦖNu�wo998,����8R����R��A��NY��W՚��JMf���*s�+u���N\��t8��CU����K�"X��_�'�_O����
:w��[C�����jj���6�q���>��ѣ������&Z��/����h}<��.S��_���<�.SM���+#W�5�(^i�|�!�epxu�7���tW8��
�ؽ}FlJ8T�F���	��P���_�c���ڇ�K�²޴�^5'�{��t���9�8W�6��˼W���*��Չ���,c:��Kz��~�+,XNw���\g��ҥ�vv܏��\�E��	'���������#���
Ov=�/b�������C��G�P/D�yy�6����f�s�_��9y�i��R*W����Ho4g�Qa�^J�}����#O.y���|�{b��>�a�|���H�W�F�c2,<<�7n��8C���~C�kk�$��Mk�?�Ǐ5��NiYY�NH`�.������q�y_q�:y�x����x�yck+?��q��3�n͜ʴ����$p�76�c:�v�u�a�I�&)))J�ҩ���x�����л���>_˿�z��ϼ����9.�VǺ�Y�Y�_f*�2L�rv�sE~�'c��3�7��溺VJ����<rD��T��e���8�^|��(�r�r�?Wy����l�4P�y����W��~�����kEm���+!�(��]�~��_	z���x_X!�:'��4�Mj������L��&��WW���ӊ*^ӎ
R�d^�F&��h��d��W-�Ȣ"�����v}�XȝH�}k 
������	���ym~��%�����Ӥ�xi�]8.3ˮ7���o�|�eF�6��~L5O�^��z�M�<o_������sӻ����E#��)k%��1���[N���h���V�'�r��eW?�{8/��j�^�����A̭�޲5����WKN�_5�&$44G!��4������<�o�E�8l�0u�f�pb�}��ʎ�f����<�1@�X�����/���PFf㩗pcv[�%�1�~�8�]n��o3����2N^)2�����(�E��ͳ�h��+E��`|����s�bfU�.�u5F�8}&�b~�R��vʽ4	��W��N?)��Ѯ�"��������j�"�E6�
t�)C+�k���əs����J������ U3	��cD���Y���Ƹ�zh����g�t�5/ru�,��ja��t�d�Oke,�m�������Ŕ���k�t(W^�"�O����ʚ�"P�=����D�Dw���ݻ��G��ĕ*�M�O0<55��'�ʕfv$��*FF/fߪ�M.u�u2�}����e�YS��7g*��Dhii�ʏ�{	�V�K�o
�Δ-������	���Ń�ߊ�=N(3�O�_ޚu��ܜ9|�־+������e���̅��1�'�.kVs�x�͗����$&6XΟ��8TB#�8:���YXJ��k�Q�l�E�ɭ����90<|||��A�pq��*O(c��-qΟ�K�_�0nU�r�rN]mhhhDttۛ;m�U6!�r�)��겑�Z=��@u�����+���m��t�ͯM^�,���pV�`#���k�"2�h��l�'��b���lzU�w������«K��^T�.|�\m~7ʚ�"!m�R�d��pHx��S���m����M��6 �c��8X


��W>���y<w"���rWQAZ��2���%G+�H�ް�C�P�9=\a��0�Y�Ɓ~�,lHhݿ�N��~�X���F�]���T�2y�ū�I�t(Ӱ�^?��g}+`�s&�u�ܢ����d?��<�|al��b="{�"�2y�T��&��^y�lϱ��#�O��{���unQczzzWy#�J�ӷF����VmL�,k]�Kjnb���'��
�X~!
�(��kQw��r�N�Ыa�u����S�OxVo�Ɲ�%1;J+��T;����]�����%��?����.P�+F������;4Hh�l�)_��S���UT�Q�/�"���t#�"�%���Rҍ !�t#�  (J��� ��-�%]��p��w�wg����c_|\0��'֚�+�Ss�TW5���q��T�n�Me\�����<&Ù�,�����4�M\Ӹ���|:�ﱬ����(J�����E^��BCCܸ�axu*���ɒ��9�!��@�����_�X�i�����\޾�̟�~��q`W��Y����C�1| �f�4#��l��vڙ�
�~���QM�467�Etb�Tڢ���gW#�֮v��a���^�%a�o�F��X]���Ctllr�����EUNp��1M-���B\��Ow�mQ�e�c��d�}�6u�5K��TSB��2�����|e0�Y]��;��3�h�`��%��'#3�݀[.Bђ��D/�I�1��lB*Du�h;#���K=��uF�V~��!~��1
�"���;B���Cu�O��}㚪1'�z���;������������h�z�znGJ����:�����\xK�;1���x�� 	ppq�'o`Ԣ|�&���EY��i[[9���1M6�]u���ч=�g�.�ca"�ׯ|�\}}�0��Bgĺ+��Fy��_Eou���p�dFټB7m��'�[��f��Z~a
���dٻk�m��Ӆ�NK2q���U昒���&��ŭ�&�|�I��l$+�.o��-�E���՚Ư�`/$��c�g�O�Qh
 �1�ϟ>}u��벸t�S9u��}r 	��p���Bd	�
�����	6NN�\L�e���"�ɐ Rf'%��o��CS�F�G�ъQ�~j[�}�=������}}�A�#T@�ƺ�ţ�)>�����]�IVV��e&�l���ƥ��d".�M�䳶4���::�U�9��Չ��=��@2�C-�x�����
�'ש�vM�o��P����Fzj�Ed�����e�����]����f)ɝ>+ީ��t���\lZe�9������)|6G�v��+�ԃS�QR�(����}���A�gNd�;j:'c���Y��A��2F�O�̔�$��LЖ�mﯱ���	�0EEE��A��y畭mmu=)���{���}���62h5حSt�ud��|,�͛7SY��uK=)�ou�V'�i�޽;H`����y����W�x��"�w�ճ�����>��Lѫt�vPΝ�"j�]���2&�&�q��@i��� 
o��g��?��(M͉͢������͢���/_�|�B���	�]�^19�y�����4�`���[5��%��i��?X���@/�3��P)�xZ���BEsK��F����I��M������C��k��*�F�W�����JӴ3���e�Ӛ�N�C���qDA�㐮�؝�Q>���.=�Y��g�>.�j��Уq ~~Xo�H������q��jLJ�^v���
�+��*S�����1� ��ݽ8���0vWW-�Ľi�bx�W�5*�g:��a�;��kԌ��Tb����W��{�&1���[hg��Jto�v6@���9r_�ހ�(�L�@ǣ!��y����c9�-��~��Š�x-#0�^��O���r�h���؎��i��۫㥄�ǇG�����]6�%���&��cfo5�wx�3�ގZs,F��ŉB�M�o�,�<~ă���y���L�!����<�e;�B�%�ܵJ��0GWBAFF"^��M�M�����=�a����]�[���ښG��'�}(�_4\�}-�2N�6�ۮB��^�`�V�؋:C���5�oT.����uzNpu���>����W)�&������Z��6���Ȉ�,(�;K�b������ӝD.#��D��[�B�����y�u�ρ�2�2���U^,0(h�<Q=�!ǯ��WdL����LK߱�w��C a����UW]��ᎇ�*W�&kQb*���T�aXZ6�Zf���RS�/u�,l�v��7�c�PT_��y�&��+��!T�ɑ9�گ�m���d'�|��} D4��a9���U��-\}8T}ިy��R.�����:�o�3�.R���D�xb��ܤ�,����K�r��n�Y��'������Eɐ�Ȳkda�ǰ��Ͳ��HK ��( ��߆�������..����fd�?[#o7�٫�ϟ?���5~��MZ���z�:��.Q�]E�������'�I�;]�c�p����e�ZЈ	�&1*�p�V�BL�'������\wnrsߨw5�w�qe�q�֏�%g��2��ٱ���B���ܒD ��0��K>}����7 ��iׅm]z^@ � ~��ugASi�ּ`�r�y�A�����f3�_
:dh)��ED�f>�����!9�Ti�Zi�Vb���z.�&<������Z�_�X�JJ�����I;8�ZuM?�\ʞهS��V�}�U�Cs�/�n� 2�%Ooɫތ��@�O�n)1�4 /������м��x�d&-�׏��v��8�0}R1ᥠD�a���|��!���|�ܗ:[�ٷ��G���W�*M��R�(ޗ7�Z��;>T�)w��]dY�w C��dDS�����#77��P��CȞ���	p�&I�^5�2}�� �e��+�)�L�!m���z٪��{��F�g��ŕ@E>�4[��O�������ʬ�W	;�eꜪ�	�h_Ʉ[E�Iu_����)���N�[OV@
_�v#NM�J��S3��Qii�y��ͦ�� ��6�����棹F�?C**D"�{�Y�#���(�k�I���ol!�� Zԝ��׏�6�g-��J����f��ю�h�W��k��%���*'�N��~VUy�^l�@Ӟ�U��ԝ&��e2��O��=I�Q~�&��t��uQ"�$YBTT���QL� -�kT�~��"2�(�$���C��y���:���>�[������̞jood�q��N����U����kA ��2� n�D\���Yuˈ���M��9���C��"����ހ�7*���(��D(��U�ײ8����%���@<IC>C��g'`�)��N�V��kVڗ���m���������̦v�t��8:�GV�r��Y�퐑����c=!��%w~G\��>c؀ê]��}~��
8ɡߔg��鰤��j���t��LVK�"�c[6r�u�̑��n�G�*\5��> �o����{����?�y"�BB�ǟ�>�`�efj���ͮ>���i��6��P#R�? �C�⬽���v���,[���U����beˆο�f���F!�uh5�?�l��1��5O>�T�/���̓̕<�@�uo�Ʋ���!)��U~�W�@����:��	�l�5�҆��>H�S]A�������2���z1cJݶ�2ǌ']ҪȀ���ܰ�����D�I�A�߆�����ۚ�tX~�}��@Ff�\���׾-�G��:v�Uo	�i�Ϥ-�m*�j��1*C�����ϟ?���J�u�pg�#}p^��2��X�Mv�k�n{��D?��Y
�w���|yyy��6�v�9�k�Z�ga��w�!�P�/.)�KU����X}H:k��_a�}Vd�*�L.JЎ>�������|�ʃ��~ �ę��dz�ؽ��,'��o=f*�}�`�^aDb_���3B/�������J��������w��nU�1G��/�Q9�^Ѝ�f�(4,�M:��DT¾ԇ9=��Y�~l���t^5�0������^�*��̑�/(�l=т�}X(BK ������ܶ� V�h�i���#n�����ː�b��,w�j/jd�I������B�b�id���a
��Z���/D���B&�yxO6��T��-�&/�/�P��\����\� �ꋃ"�P�mX�!������wP�r]�K�_�A[;׀_���ͧG��([h����۫1i��VF__h&COkV��S�4�I�'䝏�;�4F�9��{j<`.w�c.W�l����2��꾗WUꓭ�дM���>��aS���y���"*a��Y �$� �0�s�(��P.2<7�Yf6��Z���A�B�u�`�� ��{���		��'9�aI��Oc�wkQ��C�'c�D���wK���K)O���-J�=�0ntg����~p=|�A�ٳg,Wn��1�o�[��l�8?���^2��X��1������!!�N��oL�
^�4|9�š�ݽ�7q��V�x�T
jq��z��"oL�a�;o���;Pג��3!�����	Z~ni�n��J�y:��ɛ˄mY��w��6����ύɔ_0j*��e|{�}$�H�����:yA�\��-'�c�!ó���a��0�"X�A�J�O�O��R+kiηGf�D�l���A	��o����Q*�
��ܷl8�냎>A����B��������S'�;�����=>�.j���b1u+����S�������v�;������Ѧ��T�χ�Bo204s?$j�H?�%��=>F�Y���u��{6n}Gj~Y#�iu8���]C��|��SYJ��º��7��6�����Gq95����u��#C�v3��׮R�֔�ͶY��O�+T��|u7^��&N]���n��d(��j+���'J6����`�r+#��:�E�Zq!��Q�V�g�ާ)��iRD��y?��� >�	
ʯ�#�ޢ���Ϋ@Ԩ�����7d4�<�R3C�9����_"��bQ&&�N��?����8x���<��w�-�ݻ��2������#���K���k��+�Nc�%��� ��z��x������>�~�AH����a�"���
Ua���)����z��o?=�Q��$fk��e�I����� p
�w^�t��zF���
)��70����It��#b����Qp�(~��eZ�Sdd��+ҍ^w��{����R*bq���n��F6Uk�ĄSw����[Y�a�b'�=g���S1b]��2���%�G��iU��D�����&ɿlAY>PQ�2aW}q~���/��W�p�k��%ϋ����7v��c�!�1����HЧ��°$***���)|�����s�<��.wbߤ#F�4l�~���O����}+{hO���R�4d����S��JW{��f9���F�C7S��֓(S��	$]h�g�pbY-��̽� ����(��Yv��`�#�ƶS�]��8Nk8'Ň��<�jCN2�UJ�G�}�W|s���4656�6[�\+��/wL)ǰ�
��׸����`�"R�7L���e��ߘ��C��n��c������4�L;�����Ŋo���N�܏�����@!�"����F�ۉ�����&b�����L�.ΚȅX����F|)hgkO��cʼ�²'3�u!:/��}���F�pFF�BR�Z�$11���j�Љ<c\T��Λ/�5�"�]	hi�s��^3��{>��Y��@#��<۬���l3�yͦb+//�����̂��bg�ʍ������N}�ng҉��R�3�ja&��ڗV �DX���"%���{�_p��ORe5�lӊW�����U��2ֻ�g�6�����8����&�B]��:^�;rßС����M8I�sBK�ͭX-b��
����-�/�Q���,[;ZL��5 �Z8�W��24���q�p>T���:����j~W�6�D��^z�,����(��!�
��w��_v^����Α�� ���Z�ѫ�o��g?���ЈrT�a
Կ���P&ψ��u���L�\��Д���-���=���r���mt�EGGG�^�����	Ma7p��+<,?��o����$�L-�N�b�<u�(�崒_�ȵ�"�����..��߯�FgQˆ��}�d��L���W%//��8T�y���(��]��^� )3����Z�ҒU�p
�?K�|uA�a�]�9���`e,Z�%���Dpa�EV.���A96�b�,H��t�B�����ǻ�_�*�Y�C��=�R�.��z)�q`Ψ���t��+�i����g�9r�~���,���u�&.	���Y���k{"%�;�t�E<�z�d&k�n�!��FR}�D���0�����O"�4���Fzؐ�@�p���pڿ�ڜ�����s,C1'�7!���q
5�bk�
�0>�����{��3^��.�B^.�O���F-�x�kEl�dW��U���<>�50C7��s{�
1�Q\FD�����4(}���؈���
"���Iiw�Z�X411��=t���X�����U�M�$��v`38����~��aIC+�
�_�i�O�wr�r�D�&{<2?�ۗN$.&�����1�_m7A�C�ݠ���R��q6??����E��V����Ld�\�շ�v:z�����jEt�>ɽz�-v���Ѻ/������������M1�\�cZq��_1�Ǹ)=�6���U!ȣ�p��S]NC��q�n��6�½v횘��H�#ʋ��L���&�eZ�E3�w���Ӿ�&�͟?rd����<~L�b��ȴR��v��N��0R��>Y�P�������=�[�$�,�~�_��1#t��AC焴��\?"���s�Uc��媂�}��������'�ܵ���Z)))iT�p�Uθ#@�gk6L���2�z�I���e�����1>>���y��pm�h7[�N�j%R�0Y���%�$�1,����Kg���zח/�"Տ��#��Q`�N��S��S��Q^
�*n[�ӂ�Ν�o�����q͍�� ��:��������(��,�t��"k���o��D��jٹf7K+�g�h�=�v��O�kZ��=N�7J�֖S���1�R@~Ktp����,����kUy!n��ӗn�-�^R��(�2�gԭ�Qs�U�LEZ�+a-�t�f1��^��V�bb�����P�x�^�qI'hw��Y���8�o��Hj�H�ه&�t��º��%<�X
��޿�Eֳ~}��\�<:�x#}@I���iZ��]��ig\�� &����A\�@�$>� �O%����'����o�/Og��B�π�aV}���;	]�Raɟm�_�i��;���d���gM'ʝ�+{�
7⥠%���D�8jg�en��		in��a��N�Aj�T#��	���u�!5k,�/_���1�Zؿ�)f��^�����(��^�zdt��7���=?u-|̈}���Eq�i�X������9L\�7�䱊IL�3�d�>N��w|����`�R@�5��'�k���� 3N����2�!�*È}C��%o[d �H�d��^�u֝�m�J�=����w�q�?4����=Cd�v�rm;Gu0�����d��	���:�&&�̪u�&vΐ��4��8(�]�
�z\�#/��ppl̋��O8��C?��n~���su��ի��� �7:����Z?o�t�g(������7a�zLmF��m�b���W���bɏ�i���'|���ʩ����O��j�X5���Ѹb@o8�>�M�a�) ��	N�]��K��)����T����`��sGL��h*21A=�eF,,��bV�-�	��������k�>��Fn��!^�;Y�w�=�L��W��>O�LMxUbRY��˺��T,�����"�h{{{�648s�nļr2�XlL�ߡ�*��*BL_�]��J��(��U2����*7��eB�neee.�q=�D�Oc�����8ܝ��0�Wg��9;��RBV�~�	����N�@�2ݽ��p����, �|����u��}vЀ
�3$���������A�_�?7��ν��㹽�˱�����"��a�Q(M#H�/42?�h��\%Đ�_�#D���4^�D��H��R�|��v����)�#�H�L�j���.u���J�ve`�~+i�=f���������}����f�N�6����c�5���p�EO�8ר�Y�1+�	��?U��$b8�K�M"/M-��C���lO�S�#�Yn���*u*x/�K�b)�4��5��v�3��1��i�q��U�����D'�MTP��Wq����A	����yqo¯��#�ۛU��+����1$]����Y/u���)[4��(E�g���.`�Sz�<�c5�fu9�p�}���K��g}z��?bJ�T�泺j�D%OH0��A����d�u��1��\��L�-��{�;Nh�H�����0u:E��ڦ��&7w�m�/s��yt8���vk#8I��%4���(�S����a27?/$�ɦQd9b�a.q�o�A�嘮��`�^�g�1!�%|�ho'�/*g�DPA�ߢn�fE�m����WkXQ�eg�S l>+�i.�՜�z<M�+�q����-�.P��b��^ߛ�E\���U�ư��U<$jx��|P��xt�9c��͈;(�����^�H	F2�2�J���]�ԅ�u�~w����I��\VM:'/��>(��$aQ�"���0�Ў/�%�~p�>2��UpS�BYH���@C��`cklg�:?ٸ���=�N�K�
^�� (I,_-��W/����H3�De|���)UTlE�ʐ๯'�>hU�Ƃ��A@M���r�����!�o����L��[��36�ܥ��2kr5��gI��+,(`�) �&��1ύ!}�����G����x���DDI%�Y��XIp_�۫^_>���!����PQQ�.:����q�k&�7w��� �:1���ټ�|�>gcm��(�AQ��1Tz�seǷ|�h�1�w�cmW�d�o�mhH�����ؾ�Gcr��a�[�#�4�M�Ws2O����:<��a�!M�wq�HQjT�nի�}���QM�.��
�� }��=t��e�]y�Hu��?�_
�E1O.;c;xW������]�����:�<?����P���b���z������b��2g��h%�Iσ��aPHE�2��	���8u�a��p��\N��>���b(�����U�gV*��Gƙ4���1��w���δ��Ï8�ܿ���0wm[��"%o��r�kw"D��AS555�5_�cP����6F)�Tq��hQ���4�ݬq����0�o�� �>Rߋ�{ְx)O���
��.���g	Zl���	׿�dF�XT�@��%�f��Q"���J#�f �o֟�cZ�u&�d�,�(--}�߂�G�!���231i[�(���g��A|�-�H&X� �b|dŅ�vgz�s2���������vJ	�4u��9!@���	�}�Nk��#ST��W|7�d��
-�-�UI"I�.��kE�[�@��Pװ�P�a!�Ǒ���j���D�2�<º�PiM�u��%�'�����������Κ�ࡲ��^�o��D0���+Ydh���y�ԄU=>o���Ğʠ"��7��&�$�XAKkTH}��p<��yT�o7i�n�t������˨	р���R�2���_+�2�m�Y���	�$��rKU�b	�Z�ؚ��rض�wj��l4*tۧD��RJ�g�����lUp ;FFƎK�.�ʆ���c ��cH�i���!�_�cε|R�Z�,b���W��#���VO�z'5�2k������O*��u�lk	�V�..%�w��,ޤgCO!�{R�2W/�ّ�˫�6���B�FI3B3�g������W0:$_��M��y��K'�=dқL؁)999ݡ�R���~x��=¹���@ۓ�t���Y�j���x��)�~�y�y���K�45|��y/4;/�=���qԌ�%����X�D"^��]q~�����S�eP�b`dڛ< [4��繳��+G	SÁ�����]�����Ɯ�w��uW./Qe���-�I5�Jp��3���\,su�%��d��!d\���cc!�6�׋x��W`4K\�4��P�toZ�t�%�kP��/V�ݐ&x�B��h��L�Ϝl{�=R�!���p|eY���|�Η�ߘ��{�Y(�.d5Hۇ&&?b��XZ�?�U��i�fU޻���7��������fg,aj`'��Dp��ۀ�L#�ֿg��S���,Q��|�)\�ztsbć���V��B8=6��P:���b��r1o"ش���4#>%$����O��e�䤽��b���c��5S��/���Ke.����##&�q� ��ā"� *�Aȩ���K#�[�R�H��*�B疸l%������q�����D(د}���-�c:����� ���0#_�Z)sR�|����^r���Ћʟ?���ߺ5�A��P�.>���@Rӛ�9�d�dĀ�}z��h���AV��/��������-��n-&z�ۍ�P��Z �_�SSt\\���.2॰)�v�A*�,�V�uz�%1v~~а���s��Sx'4�"�Ǧ�0uJ_a
		+aY���FU�z=��ʕ�**D��˝��3�I��� u	@�Z�(���T��k����]�v�a�$���C��7����FCI�[}�YGb4x*�s�dT�� �u���������mBX3�d���DGG�ϓ���Ὣcy_��\�;-���k>����UJz11;;;��x�--5�>@��ІpݑR���r�]�[�~�8�����,��5�K��r�"B��	0<��"�B���5���MQ::ԧO���T�+��<�Um���U�;�Ძ[Zd�]�d\�o�g����iA��e�}��WQ���/ �vM]z���y� ���TZ<
^�r'iE����MA���%%E�E.ꢺ7�уV޼{w?b~���v���
%���Ce+o�N�-:	ח�hd�9�j����S��<iJ��8(��]kWn6Zp�*��]aQ���ȃ3�味�;o��D%>�-�~��?�yoC
��]��K�z@)d�s�O%�����ӏ'�$���5��_p��{�(� {� y����sh�V�����CA�������Ϸ��cY�/����T�̊��R��Z"[�11g!�*�QwM����[J�OWy�+���6��ʪ���ٷ֠��y|:,�G���d5]A/��+�k�u��{m� Q�� q汎9:�
:Ӯ||=>�S���Wxf!d.���D�LA�v%���g+��Q�Q�ϼc���w�2Ӎ؍t�|||~�Q��w/å�eQ��Ϊ�����C��� '��4�H[�fI���!�`�S�R�׼�~?��ȸv�}��-��MߟD���
d�d:�_����w��_�dM��d��C��uV�vXLT"�P��"ۏ����H@���&6G8\�Є F&�G���p���҆B0��].���vm�O���2$�}g����;
�<<�?<�H�N� *���*xii�>ɠ#!�+�t�aV?��֖��./��q椥���566�2����\�,�`�oQ"����	�ȺH���%�S���ttLL8�6Z�m���Y��-�����	Z��x����eP�M�ח���^(i��1!���Pa���%�E�N����U9��۷��������\e�W��n�H+D��V}��e�3@��P��f��'�{)��h��~d�ɺ���O^���_�$��"8*ZZ2���p�����/ց�Ti� ���\���	�H���pt����׍|�/ (Hy/N=K�u���^�!%ePw��@g�E|��eta���2*\�:����Y�*4
w^*�#c��]��#ܐ?j���'!���H��x� 
^3d�\R��-.��h�`0�(�Iz���H>��h��[��Nv��?�������U���/�H(�JHUeB��,[��ӕ=3�AvO[6LE4�$��m��|֊AѤ�4��ÁNi���xKRsj�!�@u�/�{���/��WT���S��Sb�``�e��O�?����U���0߹�h�B��C�ލ��=�L�-�����.���^�b��|�3>$֌P�����}2b�P�ŭ�?VT��$Ň���}r/�0V�HI)/_���ּ�8*,��`@��Ŕ�����ë⧧s�Z��d[Z[���N�˯w�P��L^$��'�7sȄ5l��?#F���Gfg����������F�T�/� )�c�M��*� I��?��0O
��&C]�1АU��6���M�nrp�f.J}c�8W�z��~���ph�*	�[󤺎N0�ӫ182�L駔�0_�Kb_�@�>��E�]!�Ȝ�D���F�F��
U�����ĝm��A�wCe����������p�<��i��B�uF,D���))3J8���C��6�#��*zC8�-K��t'�2Ι333c�Z�$Nr�_ӯ�d��9?�m���?f�H��:?v8!)���#?g*���/�s���:Exa�z��-Φ��U�s*J�fH�Wf���\%x�L;#'ӡ"pHLL<r��֢�C�{*�u��w_d� ���+[�p1��>�o[9�6J�@�IJ�C۟�b
��d��0����������.�Sd�$����Қ]x���Drد�n���"��w��NՂ^�7~6pd�H�M��r�+�f����Y��99o����� c��($�����d;��A�����w�B�ņ�^���ϕ��c�C�.�	9��-��wf
^ܟ'�|/��������~n��12r1�k�d�U�b0<<"��1�u�B)"1q��"��.R3hׅ�Ƨ�\I��>�Du�(D&_6� �z����q	O�6׷H����׍��&�$&^��:7h����E�9�J^J�xi�R@��V���Z�g8�ȍ ��T��Lee�Os���6Vۋ��<9����d�_������HZ�&g�����c��pW}��1-�A�'�n�E?�W�esJ�Tm���3��=�����<����zx�L3��k^���;��q��mx�"+������?�,���~�gJ�e�p�t}:�)0JؑY����L�[��=W\� �o޼%��_渲��Le ]���h!���"
��������mΣ΍�pⷤz�2��>@[�D)��6[�D�S��3��l#� [����WT��|�����#�T�/���
ߤ�"pE��~�R�$wQ�@��b�PL\��	��x/Bз/�8���ܸ��:^�qیڼge/�3��@�|�0\�;P#G��4���@M����#9����9U���g�͇�#[��!|��k;;.�{��.t�#�o�#�;�����GF�/�e��&Ë�YTc�w�Ѻr�}����3ԡ��ݻ���g���K�E��}�ާe����cd�����WG>cHEQ_�u�xw����{����8!{^g9䮑�f�ՙ�|�߷�/_\ʈ�s�qI�YaT�u5J�� ���c���@��Ј�U�h -kR@@MU���FϲC�5,D�����l�?��]�Lp�' �l�W�ɕ���D���!�� ����No�;;��)��N��2��7��sUS�ګ�����������W��qd�{~ve03�\lYn�EX��H+B��e�Ydw�������B<O����tEq�J���ش�����6
��E55�wz�::T�� e��� m���"B�����t:�����-~~PBe�I}CJNNE�h�����Y{p��&�;
�n�Nk�����&d#�S��2*�F3ȊMR'���� V|.8"W9�"��t�������v��4'16P��'�<UE�'�ϼ���k��G��4�ܮ��>!Mֱ�X9Ę�/�JgQ�J{��ҀCH��-�|?Z��Rm�'L00b����׏~�E�wt�BW��״.�s��Ǯ��\w��KJ�7���Ҙ�����"ڲ뉔����"�����\9�J��58��`.��P?������/m~�Y�Ιn���Sމ��K��KE�<&,B��<*Hӫt��������ř�����9�d䠘5�]��5����]�~�ODu�T�@�����o��T�0���L�ߘ��7��J�*w\��S��܋]�����\��1t\ả���B}o]��ռRaW#gA�������g2ۑ~�vuF^���74 ���P����������/�u�e�(��01���e~Oh�wf����pk�7/PLԞ��G��(
	~��u��PtI�(���6
�z}�@�D�/a�o��~�_���׾�3�uXܱs���)j��!f��A���r"Dd�ȅ�#��]�%��}}}���F��ύ�b��������N�_���(+�(*fm�xn�"����ڼR��Q��5���d1qq}}}����1�������������I��w��ƖOX���N�0�y��,`��"R�M������V�
$2��	'�(Yiy�����PK   sRWZWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   sRWZ��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   sRWZ$���� �� /   images/669aa2f4-fbbf-424d-aa05-a9f27f46a07b.png "@ݿ�PNG

   IHDR  �   �   M��   	pHYs       O%��  ��IDATx���y���u�����޻�{�g`��N$������T������UR��,�N�X�È�T)Q��P�rLR$A� �3�`��[���߷/��s{T���*��z�����w�g��s�9������<9Τ���D�7�l`�cK����7�S��@�M�\�~�^�q�e�iDQ�Y]��Jv�Ȓ��j:���n���fپ�R��ӈ~/g��롔A 9�ͤXUՂb�*���}��1E��d��aU?�eU�/�_����ql�_RM�W�Z9���mۆ�%I�*~�(�eY�d��}IM0��x�#��C�f
.�$�?�{�84�$�]4M���,	��/cZD�	Q@�`Z�X��/��pwU���[�G����/�(��I�cE����1����bQ�T��Vm��w#�=R�;d�2�����s��R"�޻~�R���u�J����^�Iec��>�ek�CϣI�ӄ�N�WS���h�0��0�� ���kjD�T|#�:�IR�ְ��ph�L|��=\%+	hFt-݂�Ｂ(�����Ȫ$㛼]���ȣ-�Y�& ��
#\��ƪje�S5�"�D��1i�_�\� <[	�Ǝa�������b7���e9��q,&F�fҝω����@��?%���Oh�����h�;S��U�����YL#$�E+e�OÀ�N�}�ǥ�f��v{s�,���iQ�B;"Ә 	��8GIhn����#��*��1�c��}�c�<v�Na�{A� ˱$㾊n�^$$;��j���U�ܥ��E̯���J)i�I�������zo=5!Tl"fY�HN��e���B=)�#�%�9Pf9R5|/�Ke�!8G|�Pe�¬d%��B��L�<����r��9�a�V'.�I�Ϩ�.n��2�B!���"f#�<%)y���UVH�f�=�i������e�f��*��F�JՄz�in�JBʬ
�oI��.a�Hk����`�����k�O�8w�[,C0�G����0�"���$��r���5t� ��2::
�q��u�@
}9� Ֆ���/J���hcҀԺ��`�H	H ns<)t~�.$�s��L��Cf5��+<���j�F���f�
����'f�3��)��QL� �,͙&FQ$�4'T?�a$��_��	%��SV�O|�s��"�=�/���c��L�!2�\�
2,��ɬF3������M��H1e$0X>�
IER#ќ3��J��/tk�(���5�eۥ4>6�T*�G����q��m�O���QՏT8��gQ�⥩L���B��i�7 c�
~�ag�`��იۏ�~�r<��!)�KӾ�z�B�����=�#~�i7e�������. _Ꮍ8ac$@�~��0�:),( p�4��a��a�h-����Mwgz���1�I2{h��U6ך���Dǜ�@����#�$$Cn8:n]�ڞԍf�@�8$�����=���
���1:*�VSR�P��_?�����c�4rDk�_#��$��=bc-�� ���e�~,e;v�0u��Hظ�1C�'�+J%PL���<�����gۗ4�e��l�����O+M�꧙HD�a�%��1r���.'q811�^X���S	�rF&٤���o������A�&fM�_P���ȞJd\M�d-N��1 �E��Pp��FS���v"�;�s��Bf�s�N�)��Q�PkN���2���ڠj��[�"h��N�c��{�~R�q���nI�'Ї�}�tCuSc�I����7���3 ���y�n���U?�J.�uRx�F
�h7·�r��K ��
y��qT��[iE�&�"���Leb��i��K�лGvM]�v-�s ܀5l��;�C�C��K�֔,�g����EeN�ƋYdk�P�&f��&�aC��G�^"�NX�3/I]�e09�l���d�
�H����2Y�@^[[S-�2R����4I�|���Cf���D�4���E2,&�n���.,�
SZ]�Y�Vu�.�*�^�e�����C�њU��d�� ��qJY` 7����^@�^&��q�(�X)`��������m�P�	�����hX��R(_U6��/mmmy��q�>���^ੑ�LefD&k๺���qt�8�� ���a�e�pH�ȑ7����>���ό
�g9'�X'ό8\̐��E�U��at ȚdI��d�9Rj8���$��T��~�!��I�YŨ�D#�: �d�@)g�Q�$3�C�����E����EU7+�Z�wd$&�/����Q :+)%�:S,�����K�D�4uPC�	����~�PtX+9IChUf7Il�d���j@�2fY�jK��j��|���ŕec���jNI���H��4��T\��´%�u6��|��ݵ%OR����s�ޠV.����	aհu�LTT%Ī�g9��4ᤨ�Z���~���e�&��}��b,�aG��/� ��e��2��<�9Gr��~QWݡ�t�\ʹ9A�������:8�]h��~��n��R�F�M}���'��q$���R��1�G�g�>��\R(��-������褬��D!�N�A{�w|���Zo�r/c�iR� S�^Z�K+�XLD�Bf��؀�$᝼�B��J
��R/���&S7���y(B��D��<�A�C����l���a���=9:�iA�3{�y�3>>�� )\�~�t���˗/��>@�Jk@�8y/��"D����FBr�:�H ����APRR5L	��\E�g?�q//�Hq�C�Q��?t��8R���aL8K�T$ht`
#g�G.�q&��C'�Si�H_��+�w] Ű���0z ��K�(�wC�[(��6�e#!3�QLA'�+��orI�z}�*(Ф*L�)���n����}f^��R&\�n<�Hx𜆭6�����9F��B��
k���H����i�4v�3��MRZ;T����&,~\����$���=9v�ɔ�&1�w0daPȬ��/"9c��P[�l��u�!�xF�ɶz%ԙ�P�$_"�����w�D�U��u��mb��8���?���=�m�/3�t#��Aa�McJ{�$���w��~�ڌ����T���b�A*��� ^�̪&�H�Ǔɡ�/MJ�Y(���$�"8�����9$k�P��"�1�	K��2����:v�eH��Y�@l���Y��_���~��n///�xf4[����v1��4�����ynv�СC����T����aR�v��xu�\�yiqq�l?���%�A��Iм`�A׻�	}~ꩠ���wq)a�N������i|py�i
f*d!b�DU��؆��?,��h����^ZƁ_+M�`N� ��F����������<�5P]
n��}P���aF#�m��ccc�E��lTfff�<�E䧘p{��q�^!�RU��fF��c�~�B��H�Ac}`�,Hc��6䴙w���Lop���d3JF�kk��xsN"`����,-/?0?u��U�>�&&7�ޤ���p��U�hK(��E��C�4�l�	
��1rytB�c��f��$�5
�@R��`iD���!.�>���+�A.jlnl��`m�7��R������\�*�>�{�eo�����A��,3�4�_�tSl�jwp���7]�W,T�����Y�W�T��,P<驙�K)nlI�"��ȍ7��=�õ��?X[�T���/�3���X��.��:n!wbI�d[k��jj�ܨ0�Rܿ=4 ��BF��أ~�רV��!q<�!Y�T�q��HYls4V�0txM�{��a8�?���;���ƨ�C����I{�ʨMɈ�Z&�ڵ��J�ȓ��M�l�"`�ߏ�`}AӀ�d���S�=�A͈���l���4���6h����fsv���%�U$vccsq3��6+y�d��@�
�|��{[�,�h�!�lg�m�*[K��?�BC�烒X�rs8$�[�+Jn��e�.k��
f%#�!h��F5`�Đu'�
E�����n��jв��l|9&
��l��m�L�A �䀪� j��|�L�nt�`]��0h��_�v�M���A������}P���4�s��<o���Zxf�be����.��� �*(\�����o�*{�鬎5ecO�Au�!B���C�����E�$�ߎ莰��4CiV��t����+ B�l]5Ő}��NLÀasJaI�AgH^�.vI��Ź�1�#� ����,L��%�70	�uW<�  ��9]���^o�{kY�JUx3𻺋�.��>x��+�41h1A��Ert�X]�Ç&��0���»aWD�������'o�..��{.F['�N�
u
_J?�(ee�����z����[`D�n�{�{�}�ptUsh��O����+G���/�LL�`��� �ّ�(~P@q�!�ƛc;�)�%�͌bB�+�+++kkh*�177 �\�-�C[�%6�|R�F1)��5�Ǜ���6�*�}0�p����i-��C��"ı������~,�].��Ӭ�p̡ 9�R8�o�>�a�3|)P2�)G�8C 6Rd�i��(�%�*�
��d֨�����Ǎ��̙3�o-ad���(6G�*a��C"�SvM�y3�<7771���\���>��q��Ν{�ݓ��T�7���=�H�M�N'�)v#��l��F'''e
��S
\]X�t��w)��z$�/�8�:��;+2������p���Fh̄<�B�F�t�\�r}m]���H��8�CN����1�!� �caջ��w��9=9N��b�X8L����^.T����+�To��,>q��9t�y>��@h�^,@.v��a�j��sXn��^���j�qr�(�t���|���)����4T�::2���y:�c��Z��	�v�]����r���I�#�?BUI�R��,���w�NU!�B	���ob���x�wj�;xwtx���|8(po�'.��E��s�Vq_L	3oT+SSS�c����������X�p�b�4URVPB���2���-J��%��!���(h0��щ�Rt0��7�}�ݛ�[�����(�#����T������(�U�60�y�"���=������k��6�7���36�)�}*�J�"`�� ��,<0���Zqz�	�v�
(��=x���nml��t�Y�=]��L�^U8�H�1�bW	{�w
��������iX�Z�V�@s��_�	�͆t&�@�~l�/���J�xw�Q��2,���/\��u�]9�-/�%�4�w������q 1)��~WR��^�a��G�;5����sI��}>�%�&tԦQ0ZN}J׉{�*[��ӻ�H=M���a������K�C� M�d@�
���'��(����͘�ώ��Fa~�	U26ބD��h�B�i*�x�7���/;}[�p(#QH��L�Ӏ3�Q�z03J�r��qV@Al��G�������/-�*4g2En����H���T�'��i/KÒ�MN���i4�K-/ނ6ԝ���d�8?u��W�z����yn�NQ�$#<��WHy�D�XIZ�8���̝��}��q�$!�%#�+��H�v����z�Oa�^?��٘�Zѝ2�Fo������Ų":���:`��ӓ`e��FQ��j�9:���5��_������(/����C1`���왩���S���1	�Z�!b2�X)@a)N�������ǱZ+��	�QȆ9�}`N<P���)�I�張�N#�s`�2��!��b�]��yu�t�~�k_;y�"T�d���D�g!G���Sr&��L����A�X��3F�5�+��V��a�׵b��s���`;u&PQl��X�G�5��UH9N�ؕ)�K����$�&ȣ������C����7ߔ#:��~!��G"(����ʎaJN��󵈰�x%?99�cl��S#�mE��`s��Y�>r�cG+�����C�ꚪ+V}ddkB�׋ef0�}�T�\%=Ԕ���{���{��i[���` o�3Z�w�O>��ڽ����[�N�J,�Yw9Ҩ��W3� ��(�e[+�����;��O|�lj����BA7�v��������@����0�d��Q>�J��8<"���N�ӈ:`ʉJs�71՟�
L�N\͛�*�ӵ��EK��J{5��ؑ�ș�����{R���K�]�yl��Ў����WFs0!�`�n*�F�/|���'N|��7WWWS�J�9n��R�0D��g��a��E�V��A��5��9��'���i��{0�}�EqD���L�,���dsX!�����L��Y���P?�:Ԇ���	+ETC��c���]�������O|2i�L����_��?��?]oSLY�  :��\��#ssӇ֣���2Bt#
h���������ͳW�ST�6HӸ>�|��SU8�M�[�Y-�흞�<��v.��ƻ��_�X�����)���L��rh�q���lN�Dd�dUabX��ݻ+�&�>����������k�<���{\�N	��E���	��'Z�X~A�CSS�Vs��0��4�ՙ7�?���a��Ӝ�D����*T�̧�	��¹��R�u|p??��ը�P�IF��0��������|f�ǎKQ�����s�d�P!} 0���,f۰M��BAǍƧg���k����Tw0���O|�_\�����B�y@��P3�JκI�=�qv���97���A�c8������;��~*��p_�)ҵe�Y�U���Q�N��6v��9x�%��LM�7����`Y���̧?����^|��ly��n{f;��Q*� ꁤ��w���)
�vzPʘ^�^���z����H�����t<,b����#}�(L�)|r�&��jU�������4��֔ft���BIA�������F�5NgHfE�>��;/K�Z�w���'�eL�����z��i`��������F�?�!eO:N�M(H; �?p}>���<�1�?���|hvǁ ��S0�pV@�����gϖj#{��y��
�p��*e�e����vRF�T��)\�q�������G0����p&�qb˸y�f�� y��'?����o^�n�f"v���0(�@dX����ێ*�b�Oks��t����=r�H�h'O�ľ�ω���T���4>��*x x��~L^�h7�A(Ne�O�S���Ԯ��������x���<v��N���8�^++���>��H�J�!�8[T�s8�s"��W��w�i���ڥ��7A��U��|Kw�3��v���y�֕K��ђ�__�Q/�����7=5�F"�`H��J-	/���r�݇��_��k��%�lk���P�,Wee��.Yն?��C`�v{	�wz4�9���)�0�ު��7>������1�Z
"���i�K����5l�L
��}�櫦2���C��y�;u� J���.]�4Q-<������dN���^ΪN	�ت�"��睩f���{�tؠ5777?;��''6�~������<�������o_n�̬o��BA�l�Jhb-��dT���%�;47��9���܉��kU�Li60�ʽϝ;w���?��/�o$�*
N��������1 ��-g��
LW��=���||��cG?���{J�R�T���R���b�V�Cg������W^у��me�'o��7E��w��<t����?��$O;277�k���E���i�f.�X����y��~��?��O�
z�~�=�*o�Xp�Q��4�E-��scE���ټu�T�{����Y��w�Gˏ��ʭU�]�P���G:�>DT"G?M�vn�=Hl�_@By���=ِ׎��c;�RŤ8J��7��߽r��>ս~�ĕ�]��=ײ�Ƃ3RD��775�ؑ����պz��	�����]���w�z��g��g���_���BQ{ժÊ��{lM���NY��f'��v�{�fև�\-`��&�
#:A�Yi��X:����G�~�Jl�N���N҈���i�I�1��S��c��7�P�����9ҨXPU�2a=z�ݗ/_�x�8�g?�n�?yy}�����x�b�1�|��{ґ�j1w����Z���c��JЫ ���U-��Սa�N��|��[��̳�%���?lnTf��I;.y�2ח��_�K�Ξ{��{��������p�ܨ@*�4������?��<�/���}�{q
WcPiNᯊfSJ�ץ�`kFi� SwO �ɣ�t���W#�Șua�Ξ6Vʆ�?|�S����׶��V�4�t�S���<EM����X�T)ܿkzjd��64emb�#�w��p���K]=����q[O�K��z[�aB�9[�EMaC���31�\[[�����Y�i�p�l�Y�'�	�1��k�m��Ǽ���g'�;��d�������_���!�G��r��-��z�ip�G�Q�3 �|��L�oW:�dJ �z�����c*;�V�2����Y`�C���R@~�L+�M�0�~@e:[r� | ;q������Rr��]A�mC�$�zc�[����ӄ��܇�n��7E�M (�z�- ��{��N��p�9��"
�ks���8%x'"���f�d������O����>��O�|�<��z�Xd�*����q,(2�2(Y���H��Љ����04J��Y�'�}fR��u�ƍ^�OǶe
�`bM��Q2�H�/Ifff6.�	���&�Fh����'08=5)&fh��Ї��헠nn�!Iw�E4"J�&y:�gg�v���
�jP�FFy��&����ąE��SO=�ꫯ�y:H,Up�f�w���K���� >`����*�ya䇅B�����M����:����0S�]�T�Epn�k���Q����G��ۙ���w���ӶD���(��A
���O?���Ϳ[�:�{@G���m�ӆ�ܷou
�C�=K�X�G��}��۞���1=g4#����ˢ�� �'_j����rvf8����fBר�]����>���0�g/_'�H�����v�s����]�����9�]+:�K�� b�ݻ׍�w�y�l�?�я��7^��k����K#`,A�\��b��.�U(,+�Piޮ�R���{����W�n��_�%��c��!x`l�r.(����h���O>IY���UM\�D�)�_WePR&Ǩv�\�v���ţ��bu7��[%q���-p!�ơ�;!/�%�s�A,-礞�(��RﺹՁQQ>Ǳ/����?6�w؀@���a���Z�DΦ�P��N�=|��狵w�}�ͮ����/���*r)i'��`�i`������sp7���IՒ8n�Ͼ,M5@:�ȍ�M�c�~Q��큑���D��(�\]�6��T/\�0���S;���c�bqɃD�H2�3�5	�X@�����]{gf�dz�Xv7N��W'�������\��c�MN_c�Z����4?��F͐5�\�U	hY�{����]9{�����h������ �:|�(�ti�R������۵c�*9�t���|,��c�J&�T������/�rB
8�t6ƅX,l�eX��&�vL�M�4n�{4�938@���D�4u��*�!'��j����/��R^/%a�8W��'M�,�dp)R%��i��k�י9�onfRIC��t��D�E��ٱz��F����Wc�(�����A±���d�2*����;�J�t����Z�68��O�I�%�r���'���ͫ��w߽�����Hv�d8u�B�H��0���QG��#5)	,'��H	!�4�Y.����&������/����J��쫜&K�Id���3Y�����]3���J���ȉJ�:0�XI��S�#�����e?r���~x�T�$�29|$�͓��Ve��]͊���<$�b����{cw�L�D���C��?��}�¡F�%�݂Ӣ�Sl)yfF&��AYY�v�����޽�z�P�)w��3k8��7��\R)�r�Xkm�G���[Y����h�:,=���v=?���3Z+�??;ZtJ�:ެi��k��p8���٧���S�F��?p���3��i��|��Q$Z6U+L�(��!��Lun�q���JѤ����4�����7��7[WVn�9�,;�7.K�#��^%Q����b�������n����Y�6-���d.#�DM��WJ����TJ?x��������G��3W�B��I7a�8� ��I%뮬ƫ��F6�ha�������`f�(��G�6���#���w����wu����w�=}Ev==�d?����(��tti(��Hs�zӰ��R5r虠y6�%��B�����koy�����g�¼F�x>X�� !4�&�պD5ǘ�98;1??cP=<���x�vL�����9U����`���N��փ(�z�ՠJLHX��h����e���ｻ�ө��a4�V�Uǎ���� LUB��_�����|��^.^X]�����W �l�ӝK�`Y'؉oDf��E*�1�; }
W�I�r$��K o��v�������Ұ��M��_���Ñ5�Q^�H,�ض�!���t��^Z�FQ�()��m�'�= P4�S���B�	G� �'��C�>IXέ��Fv
�2ޏEQ�B1Dդ|���e�A�WX`�LL/-X�҄hb:��33�ǎ<<~�8��|�
Pd��<Mg�1�����a��{���P-�D�(�'�Ҋyj��	�qma��<U9�<"*��4��^XզB� =�����,`մ� �aA(�O.
��ŷA8p~%��ش�y�Fx�"`�fgg��((؆�K�&|-F;z�(�GZC��T�Q�f�w9�-��i�L������0p4�u{='��=M#�vZ
8�8v,z�����^~K��7�� ���˙�^����4����PY��cDj�\ v��w��m��gte�*��K�n{��}p)�E�:��A�~r���cI~ 1KcX��E0��3g�<�4p��[�"	��R%�
P�^���8^��,u}[�]�%hݵk@���*�eV��M���U�R]��A�r��-���%E�]����NQCU+�"@��}f�`���i���Z_��5�����uPu��9��~�=�,Rq"�;�4�0�B��3�<��)ᗮQ�d�#�|�����2ET���>
�Mm����Q�)�S`%Nߒ��i��y�iL�U:�N�4�s�G��"��B�UQ�@i���IfS6�@L*a J&΃�_y�(�v��!�~�c	q�B�8�!�Z�,;��a���v�R&4"��C�:��_�t	J��������p�(?ȭ�$�^�1ַ��E���HA����T���'�VV sl�/��ۥ7\�&�R ����%�GJ�+P�e^��M�T`Fՠ> ���(���Qp39R��A����R-!e)�adFԪa�>j�f�ݚx��r�J�=?3������l�������BM���<�(���s�����]���P�J�`Z����)�1��P�Z:1�S�m��WF�Q�l�24�i�~ ��� ��h�l@:��JN�-�V,ga<Ҭ��V�A�!�c�`�X�T��m֫g����nH�ɫ�q��&����X(ԙ���o_�����03��l�3��
����?u����c�q&O�?�PS!r�4����Yq�r�RGY��CUm�tj$K�$!0f��m%TNi7�^�]-� ��\&�.��*[ ���Sh(�����r���Y�)lrH8�%�:hE-�f�#��f�x�V�P-υ�)0�^�^��'%�P�h���;�����)���R������#�굲sk�st>݋���v����P	�����FM%�l���C�ȩ'L2j�@6R���_-ۍf)��#G�y�o�YQ����XE�4&������H�D˩>�ǂE�o�B/ʗ���B,�J�p~f���+0��-�/�����-i����?V���7̩i+_`�@$.��W�8���"�$}��̩���R���E��$%*xK�q3ߓHK�"�7+���Su���*&�k
���׍$��N�����v�}���c/��C��t�{D�݊��z�'O|��������kW���
<O�J&GS��V��k��z�:?�3?:Z��ƨ�� �@M#K��4���^d��,��a��h온JJZ)Ŋ�) 
^�v]�25N�:?6�+�DJ��3�>]�+�B�Ԉ/���
�?5v��&�d�a���Jݠ�QT!��TK���v�ӣ���$�l]SS,�R�b��h8�"�7��p�dD�o_�\��f@��T��r���D��;N��O����u݁�xa�ߜ�ͩ��%
%1���I��I)a����|�F��F�iZ��啼#9�X���`~�o�Ugp� ��Z��6���Y��>G2��\��*�R4n�AR�?3�0�w�:�̕�)�HI8���E��`綅��x�0�b	�%MQp(ql���2:�S�X�(�9є�.�Dm'�#f"z��LT�+H��L�p����޶�q'�XV�-���p12����
��N�f��E:�.�TU����(��+�߷����ҫ�`9����б�����n!�C��i������O��4���L���>|i�a���T�Y��g9D%�6��aq��a����X�v0�vX�D|m�r�ena�"gF�zc-q�#z1~�8��\1��D8���&`�Dķ�;w�y�PH�AxHP7�����l;ǆ�c�_L��w{�/_�9M��O� I��{Q��A�ߺuk~~^�-ҸB��t��l�}'�Q�:f]�1i{��r&���i
���	�>��mn'���LIB�E�L���%���R���o �Y�0��\h�R��yqd��w�(���R�fDN[����%СT�ŬZm�vY@<��_̕��\�RsMJ� 	`�x��X�$��F-_t7���H�ȸ�K8�D�	C�L��:x�Zݳ��.�j���0G�Z�mE'�zB�й�x����pX����k�|�6���wH�[4��b�v��A
"��������G'.x-X��B����RB6�T�~Q�Nn�gY*:Gqߠ��9:u�"�vu�7y� iT��/���>q��4!e#�Ts	���8E�䉽��a���JI�f*;�$�����0:tnD�J�||:	)]z;d�lGZ��R��v���S��3��r���~�(I��B�N�u�:W�2�T:O��w�;n��Mu�\����L�"�Q�0(�RE�e�����]ZY.�K	L�rj�,(v}�؉>�l�67(W$�M�c�Fz9�Oh�ϕ��?��
hM�������,3�{�ʉLn����D&�׊֠�C@>��\)E�Y��9\m*����"?��nY7Bj������i쑓��ʰ�� ��u[��C�Bj`��&�L�$�kYO�:\��Z�P�S�E�h��mS)�/W*���W�Z�j�i�k��	���aͶs��<�l���z��7
^���qE1�@o�?RU�V����Â�CN������'%$��&g������}*��X{B�BG���%�������Ā�b�.�Z�^\˝БO����)�'q�1��k���F��OdЩ8����L��(D�a����&Z�$"��@J�^t8���*S�U*��W�\�yŮ�Qhiz��b��d�*TK�¥F����P5��
1u
H%=��kR��Q�F���hc��K��$a1,v|7�n�����X�p�������)>BT��
�ɐ2xZ����?�9g���Ɓ+nY�Z��S~�Tnd15hJC]0׀>r��j�k�.���S=Gl��\� ��>v7��)pzt>̼y�o��b�XjG�xC]�JE�R�(脫N�V�tq�&ܗÇ'��b��M�,sgX�J����olf�� �y��I�A�S�������` iv�� 
���az\�j��J��5���.��k�4�j.u�2�����Aw,`1�b�*���v��/�J�)
w\Շ�~Y�;J���M������Q�ʱ��15��:�$��!TZ�H@���[:&\ޕ2��&kH΍#)����P��#�=��`�@��f;���FA�h��{r�J�����LxG��T�Hݦȥ�'����HD�'� JDE�$�S{E�\�r_�~�RkL����*Z�qh*�M�� �@��˙�F��Bq��R5o8�rT����L��?k�oS@�e���qY��}�ᇕ�EK��ۭ�F%�1���N�to�R���(dg8"���J(H��:[�rN�4?��BM�"?����իaB�Dc���Ni�<�;�`���<����V
l�Q�Ԕ��b��Hp;22r��	�GW�f�曾w�MMMid�K�p��7��C>W2�h��G�{XE�n�YR�Ԣ�Z�*�-���4
���LgB$MUqy�놮��~��.��|B�P'�p%�6��n�:!��­ݵ^�],��{%%.��O�.�C�*�E���37~�Y	�/�w� �kaa����B����Ab�F��)DYdPՊfk�x�ϟ�
��[["v�1��F�}P@+�*�)W�Jy�`o� ��H$q���L`J����:� %@}�g�vȋQ�+Q�C	HX�पsە
�R��y��� ��^2_P.�(�ƨ$9�Z��Lj�q����sUxɧO�؎4k�e|jEJR+����pe�|�I�/-���eH�8ha���]��~��p��e&�؏�&��M�"�Lv�!X�СC/^<u�����Rwȡ*)�Dkh#����k�p		�DꙊ)@J���Mvݰ����VV��q*�"����KU�#1U��X�]��i �-q�?�&Q8F�nܸ����Ǡvd��ۄ�r#z(;�I}B� ��A����D�/)t��aLͱE�Џ��U���3��)�e�"IJ�� �mK�8lJ��n�͍���̤���n���a�[b(Iۦ����qZ~\���]*�[�\("5ɂt\��^	���9�"q��br	?G�J��d���eml���˓;_?y��F0W�l�e�H�G����7��}���P���D,��k����6m�d�6C/��4k���l4玿�FGV6��dE�ɘ�]�����R��޺���L�.Y���S�>Ho*QI��С��2��¸d�޽�Գk����S�b$>��dTIy �K�k��H���(#ۉ�0pm�����ȶ��Rz�t��͞U��W���Y�-��;5K�"�`e��aZ(�'�#���v�,BY�
�	��82�T����j�>���K�������G���	�IM�fdJL�X� �y��O,���]]\�/)���Y���S�^,_�~���*���3��\E�H髁���&����Û��"4]�ژ�����K�;v��n}dd��̗˒߷!��1�̯.^[��s�����ඃ/���wG��	�5(�N
G&�;���W�޽s�ߕ
�)��~���RBOMX��,�|�X�؍�����Y�OD:��H��/�I@��"Ϊ�9r"�w�w�^�������[�j]�+�N�ũ&�?�[��z"���Kk�/^��Ґ�hue���'Q��j�E4Veǁ������{~[�J�*QX%AÇ��&��7��+�Μ9ssy�p::�\��� �F^ml�������{^Ώƴ>����._?�,��ɧ�n�
�=;v>���Yʕe�9eR+z�-��d�����+|��7Kc�j��{�F�Q��b@�H�����D5WV[�Vot��3Z���/����eSG9��@X��v$����+ѥ����?jh���֪�	�.�;m��Rp�bΌ����ry�l;k�sɚd���z�9*�$6T�)uLR<ꏯ�V�5A��T������1?U'�?��"R/3-�Ϥ����j6�ϝ]ܐr�|������zkc�ZF�i{k�X2M۾psu T@���=fV��ފ�Qe|�z�OKd��I��ĭū��h����k״��� �j!��S���)�w��o_\:th��FB#��T�*2� \v�?
���
��?���m�\����Bؓ#{j�Z�X��~r�Y*��Tp�0��U��۶Շ124��7������G���5I��X��^x�|�g�|�h��A�j܇]2Lɶ�R��z��������&�F��Ί?�����y1�v�Ǵ��|�c;�����u�o�yz:�\�X�$E�	���ZwiiI�Df�C�	#����Ҽm@�^{������|����bт/m�2*���f��ΉSq�b�Ƽ^��(n�,ո;��wc�/~�����Ⰱzq��S,�AT�S�����v��Y�&5��a>��������
h��>��/}3�Nxmm׎Ԫ�[�αy������=���o���µ����N7��N�z��.����Ї�8~�(���T�)�A�z�D/7��,�9 ��cp�IFS>>�~�+�XtRk}���N�<}�]{	Kb��E�U��p�k��]�v]]Zz饗t�����p�>�[�0yp>/�>����գ���A�$J��g�\��1��ak�����2�&'l�c���O=��xz�Ia_�v�Ь ���X�_�B���s�QG �ZX=_~�%�O�8��T-]��&��O?�GAY�Wؑ"����W�Bρ	C���$�NpJnǩA�&kf|��Gf�AGt@e�`�ްw��Mx���{뭷�{|	V' �ܮ���awH�jW��k/���/|�	@�JN�����s9�mG�����U`�_��_{��c�Fez�T��w�"$��Ʀ`�)D�I��2W^XXϏ�r%�b7r�(�S�[ 8�C%� yA��ǎ�fj���w�K��m= ��@=#����ɹ�dJok�8>��+Qg\,��������%������]�.��9ꃔzc���W��_@�Y�<E����WV������/����Cϰ��ޑ,с������&��a�����:�\���x�k�RJuUe�t����a�!��OT$�������T>j$�YpM�D�®�.T�T�-�}ǻ��41R�N�@�*��Ȣ��QU��y�6�к���i-��Rc#�+$|�N}Z����}jj����/ܹk߁�o>�B��5)����EYY�%������܍�n�=��KT�
6��pA��r���Y�0��W���uxǮ�W�x�V�a������j���JWV�[Ap�µK[K�?����'�{�ê�{�$V�,��������˫	`L���(�0t��$m�mO]\]щ�=hmn5l=%c"�r�~*z��u��⍥��C����ݻ�o�X<*J��l�9�w��S�΃Ԓf� $\.Y�b>��$;�N�*�a��Ϟj��y�_-��{w�h���C��z��0x�A��p������*��.���"�)eu�W��cR����g�}����8~��\Y_[��D	�3��n�Z޺z�j�:~����g�Q�CIM�������"�॒-S]�R�����7���Ǿ�կB�<|hi���mV�RH�a����tQ��=��_�\VG�P�0vԯ�����P�����^�������=V���羻c~��Xӏ���U:5)�+�Qr����*}��ف:K�YH��a���0���>
�ŝ��[������b:�O���z��P)�(�77����������N���_S%�2l� A�zD�l8����=�}��];&��z���Uk����iE@�A,��f����7�{�ԩ��bݲ� ����޵��
.����W{0�Ͻ}�W�W�sc�O�,�N7��8�q�rkq��յL.t��+�����w�؁�	�!�T�*�A�3�v��F�t������^����sc����K�<��\P�}_�M̼���7�\Q����ˌ4��7�{���`�!�6�0�c����+�
S3{�;{��w�X�6�)9ZJ�+�a(�u�Y��c��?����СVo-�#�{���:~&�d2�Q��9���7|��͜N9冡'�.�\���z�����7.\_0����l(�j]�V*9*�Q��#C�\��|��ݻc}D��S2G�R�<Ȕ��vq8(O���ܥ�ʟ���߹�խ��K�c��đukho�:y��G��7=��jW�CwH�X,;��EԢZ�P�:�������z(�O�s�ș)�»v�Y�͉߹��F�z���	�E�l�V���a$Ν���/he
K��y���3�nK�\��;��;��ۿ��SO}t�k�jܼ{��Ղͨ�O����V/]���Ab&bd��)����A�m�"n
�+Y��������g��ƚ�<�|��EL�M\��1}�0WJ8�ҥ�*)�ԞOLnۤ��ු:n���x�2~�7~�w�w�3 >5��Q����|�ry�mg}�׎?�E%���	���p�3����c%��_��_�J�O~��S�.>�����U��ǪsUj���;vlc�M�;V��&IB��� N�Q��7����_��G}���5��p]]�:���ـ����8�0:���*�:m�2�)�D�`���'���w�s��#G��j5j��ҡ΅k�)�oS��o}�e@H�
u�Xx�fP�~�7J`l���}�^�������_}���;rp��薭�oa�^@iZ�8G�}��㣣��("H�����;����5���ꯞ~��>���z�����1xjk���0�a���0�'N� ���P6������+h�A�#�D��o��o���n��`��V�����T&==M��c6l����(�J��q��i�I��R}��]H��}�ݷw�p�E]d�&۽ ��y睯}�k`���( �����")���sP5{����\��3Ϭ��֯���m��O�/���e�I�m��b~�Ʀ৖�\)q�΄���޽�x<��H�z��*��=/�z�*9D�N���WCj��EY<Ummy�z��M>����o�L~~~t�FO=�頵R.n
Y��r��������m����[v����d5`��(էf��/,�jí�]/�yR\1�� ��G�d���w�!r�+��oan�
�5ץ��\9����ɉ�.��km�ة�>���{�'�x&f��T+��%>��L�X�ʕ���7��g�5\h�>�{2⚩�g�Q�����������p����*^��P��+��8���#}ٸ��)��t]�M�|�ĉ����3�4�@�#u����J�U�8s����?NU�X.���2�$�À$��oM:����}w-�>���W��V�S�����uZ�bW&�ݒ+gW�6�>}z��Q,SiB7�"ՠ䉛�\LK؟��T60��4��_�'�?��?���2�s~eiqjznqe��˕FvA�\��|����zK��b��r2챟�S�Bj|/c���J�z�yk��x�����?����i��hR�"�.׭~��y�Cw�}���^��yJ�قQ�Sz��X� �ґuNT'{����/M�z�ч��=�$aNrN9?2!e��o;}���K�3��i�F�b�i�?���W��Z9G�f��k��>{�����o�7�45���wN�^��XıI��8��+�_���V���VW1�qc*5�	#����8�Is����_|�_��w������Ͽ�Z�_�b����nFQ�k�N?�n��b��a�V���f�FXA��J���h�����x�#���~�0����A�dy���3W�KМ�Ĝe&rK���B�39_k�#�\amk�շO�j@I}���R=Z�A-�b�p��wϜ�l/\Y�0T��L+��{�,2��� �A��4���+_��_���G�=tׁFc<v�o|��ɩ����ѭRel�s������P�5t�Y��l�p�R)4�5�T/������w.�w�'n��^|j�Z�&۫˫ .=�ěo�>���R�>I4�ǈfr*o�א��:%t���ȅ��k7W�<x S��^<qycn~?�:���ăͺxu4?yqݲʥ�9�?��6p�(�:�I�a��ƇϹB�R�텥�_=96�6�(@�¸��L]���}e+X�u�YK,�������������+wW�49iF�h�%�@�s�1`�8}6�����������5`���66��l@ @�ьF��'u���{�[Bߞ����sttzz���zý�}�{��<~����e��o�knt�xz�x�Uy�y$��mij��;w.gRJ�Q���Ɩ?<�ɮ��M�R!���x<Q.P�$����Vu/��቙|���-jz�|tp<Q1��	`�]�رc����|����E?����8�q2�Y�A�-Y�m���`�`獵Ǐ=�|�[v��5�����x��?324{��7=�<�س�Ϲ��o�6���%&��r�Xn��Onݱ��O�'>AQu�PGc djH��O)Ζ,�A�R����8��{�;\cH�ſ�^�w8�0ݙ��%)M!h�r0W`�V._1��[V({�X{8�t8�Oyy�6�,,1f:�6)�i��7�BW���p�_��G�U�2�kcks[[�?Ő�=
��?���X1-/+��L ]�Y�+ڧ~H:��8p�7�u�Y矻wq��޵k����p ��˗K���e�3����hѢ��^��c�hHD ?���X�b�"J��E���2;t�%�)1��ᯙ<��N��^��^$�c���h?���'��줊sL��r����oh����c���aU��L��2H_;���@륂Ǒ�i����wq�\�R(~̖a�F�c�����S�XY��M^��l�әN+�F�'�p��'�x��k���pt�Ϯk:���x����<��$��h���pɫ��f�r�@��%��{nW�<t���0���8>�-U1d9��[*UGH�d-N��g���.� ��q��+C��]y)��<^Y*Q�0aR���T��%���4]���:!�]��X( �D ��~�5� �b����΃d�8� �.cow�
s�by�6���,��%<K,H�LS�S�+#}0"�::�~�Ǯ�׳�>�_Ӥ{奮U�y ۩=u�c��3��$�ڃɀ�o�����U�pG@E���M6;��<:]�����c��o�B)Z:��!��t�<,<]*�wM��X�2r���;�`��+�[��y�;o��DK" :g��ݻw��;�(��4�#����t6�ou�|X�0�[�n�hM㍡��Ï-X� �0���C�r��91��0	�P�H�q}��c0\�.Q�����zC*����;�-^������r�2��/	�!*�#D�h��\���J�++�iJ�u�F��W_ݰaC�j"j�h8�~ɣcz����xa���/�5�߿��x<RY�;�g]�����[/���s��_�Ec3�|=���I�+��N���<x���z �{V�y�D��Vɺ����!�tE��z9W�r��`65���Ѿtnp潕����`�kVua��>��#����\M0]�i�I6">�������Ȣ��x\IgJ�:��o���"�<�/ҶF $�3)5!I ����X��ꘆ�;���1��Eʀz*nn��kEG����m��љ?�Q��R�HCWsC���쐍��|�Iv��-C�Y�Y՜��S��s������G7��:xx׾�d�91G��D�eG��|)��S�EM���cр$ڔ�W�Ya��s���m�eub$��҉!��ڽ�i�l!M�,e�&1�����2P�a,q9(��߰ER�rIx�X���h�Y
K�`z<ã��Ó�o��g,[��;;>��V)�Ir�|0���rU� N ;�xn��Y�O$-o�1J��lK.����>~���(�V!��j�C�m�ohj ��@�6L��V�]�қ5m���D�]��*����+��z��1@Lk�X`�Ӕ� N��JHA���X�:�"rO>����DZ�"J���W6�{�:�%=P�D�X�Q����+��?.
�(�Z�2�ϝp���g��[��JY��7��=��ڻ��x�T�`�4��ŧg��T�m��
��,���帲�o��J
�wD�,ޱ���b��]t�wfpd�ӀU۸Y�ѓ��0ߙl�����8�r�\����Y�c��hDR��+��˅B)p�t��{��]M���9<8�V��k�\�9�dG����9Lч�eŸ��DK�����ټB�o��n�p*�>t�o��ޒN����y����oq���&��];wP�X�#�������������X� �8��K���v���s���h�����jY���C�����H�į�sS��Pͪ�l�x��2jNSC�1�=^q-��eVzXU#�B��W��R6D�����'(���jMWDτ�P�Z>�G)vMt��U��
���d��ཿ�pA'��9s��t#_,���#���޽{m)�J���)<)�|��{\�1Eg��K�gV��/���+##��~�;�kk֮#�d�RA:���9�a��p]�D#i�;2��&'����{5��N)7�F��	�)�WU�s�Ŷ��S��f��'�G2jii�7��gۑd L���jgC��Z�i��EETt��30> C_�	���C;���ϗ!�qxr�KwA���a������oEBm�h!��"$N>�g�����S��I%�%��%Z[pG�i!�����"Q���[��Ε+��ٛ�(�.NT��-`��/ �oY��hQ�X��vC�s�z'}Qb.�V��Qyx�'��Y�4�N%�}��[��h�
fb^`m,���}sSw=��e�."��Q���E�a����q��DT^�z�$�R��7�u�i�P�t(��1-�"�?E�@5�������s�H�[���s�Sp;��ut��l�O�>Q�$�r�*�
q��x��0:3s($<���}�w� �8�RMMau�vK����s�h37W&e"��:j:����^�xG/�	�7�ա?Â=���hU)_���gE\�[�QY�iI��$B�\ j
������f:;��vs� #�OҢg���E��`�#OR��B��F�y5D�� �Р�ed�i$R)#���9�����ir$,��a1?յ`��Z�M1���4�S�P�b�kib����WhڤO�z\U�gA�-{_�T�K�K��U3��R�Y`�Ғ_%Lj��q�~�* ^~����c^-[��whd��f9^�3z���E�eK���-��\���`bזFɄA��ND�9���A:j��)F�x�[�l�X����+J��bgg����Va�w�9JD�d! ��C�����ªj0�pSYpi����
R<�8����N	��Pix�^&~�RΤj���
��M�E�Q��ӓ�pP�c�Ν;0������:6%nT���L�%9 `y>e�6s�G�>�l��g�y�������D�������-��Z6f�G����o�;m�S���ōmGxzlLD�#Txk��)�RK+�5��Qb���s�R-Ef�Í�e��#vP96�׹��3V����gx����5K{������4�
%l=��G��RI:jK�ZF]q��?���{�S��{!~�aej*�(�/��[o�+�BQYR`rӓw}��oGG �Q4i� O>�l�p�P�dz�5���c7t�_���}mfl�)e�����F�w���ɡ��=˧����1,�X\�?����{K�
z��?��;۶e23u��jAkhi���?(�w�q��H������]�n��J��P����͛7�#Ɇ��Y��7�*�*�Ubۗj��7�ܾ��ד��05����� ��j<��n����L6=��ػ��m��D�elk(NB( �5�g���P+�̛��ojjJY�����cR>�����YF����O�(��Bѷw�n۶�1�IˆN�$�mnd5Z��JlH~������}�3�V������0㳳�=��o�{�Yg_w�5hI"LZ���|�ٯ�¤�*[��d�Ĺ�^�#$Ĭ�׿��Φ:��K�p�w�����<
ө��睵dŪ5k֨�ċ/�����
�@�!��}�ZSa������X���Kw��֖��P�y:�~�oE��� F|����u��Y�L"������d.�VmުY�)^F��0����sn��v�-ږ�6��]��l߾���~@��io箻�
Ǣ��?G��V �s̚P5Ӡ�,��".)R�BT��֭��>�[�,��(h?���BNt֯?�o!��{��gw�=l�ɖm��X�JH�Y?�(�k���X�T����㈝9���N�a�������d��-삱�Ց��xe:;��Yt%1�
]����8�ę��u�Y������tz��a�45���NN����?�ڽw&?3���{߻������﮺��y��I�P]]2�6�~�����
��Z��o�-L��c2�����ܵk��^|~r�Y�f�����D�,`Fm޺ �߼;���U�X�hx�d��ĉ�}C��"H�_��a��%�F)�ab|����p����;z��~�ľ�ۍ\��/|�r���A�?�y'bA����7���Dhl,S���9&�>���C[��4�8!4)�I@4���=���ߕ�K��~�]������M�6���%K>��O���kc[�)�&QcY�R>�u^q��� 	��!v��'N�x��꓉c#cp-�I][ۂ�9Gz&����
f�\Fd��7<=�wC��:�)�
e��`H��S&IY3a
k��L2�;Ʊ8�)2�,�?E�B���+��Ƣ��5:dǛK�,�IL��L�x2v��z2��
�sΊ+�����GV�^��軮�$ŋT68��ԈH�kpU#�@i|wlzr˖-�(�[�-���$������(����@`��' �pɒ50����=�����^�J=��c��?��/����*������ԧ�,�!�BOO��\
L49�E� &�:�3��<��b1 :lϗ����i�[2NH��p0�w�l��^jZ����?���[:QU���q��TA�Hb�"!IFn�J�4.�᪫���/nzj���xxQ��U��e�$T�B��'��S��̺�Ę�=�*�,�8�A�qG���1:�=ܺ����#�� ���I(�9����0�Y�S"Fz��u��dD/h�cٿ��oq������G�qy�W�����̛o�I넎�N1)z0�Rl��u{rc6��?C��ц�������O����"^��f]]m� &�9̊�!�'╀w*�-��D��U5���$�m��᫯>��~N%��,8��+�8��p}��3-o��rEdx-J��
��U@.ft4��XW*�Ihε�Ŀ�˿�y�0O�]m;v�&��_���peƧ�K��`	,��e� SSi�������l2��nL=�%�\������K/��>>�h��;���_�r�~�m�B�<~_=ِH��n���z�0Uٹ������gAk��yIG�d��/~�ͷ<�"MOOڀ���[�e*��56F���'�_{��Y��N��DT���t-^ܥH<�۪U�֮]��SV/�ϱ�"z{ǉ�	3۲�Lڌ��$ϻ��A�X>���&�@+A3곙՘'��o ).�b�7���/����g>�xq�#�n�P�OSp+"pl����Ł���a-fI_��А2�bcc���(\w}}�d߉����n����.V��;�o�Ⱦ}�0�]�{n��ֵk���X�!�0���4�8�d�.ՃI��G��e�OF�]{�����љbc|׮�0�x�Lf�����瞓��w�`�����3�h��w�� ӈi�e�]���}���j(k�,�3���&QM[�#%[�5Fb�:�i�1V�H/�'��J)��G��k���0Fm�]k�9{x|l��k�.-��Ke�'�X�͍M����o���3S�道�*̍��܀%�P�8����w�?��1�.��r�[>�顑	N�?��/̏ӞfffJ�]Ep�v��t���E'��c������8��Y���ª�t��_\���9v���.knk����XѾm["���KS����h��������Ɔ��,��wO��`�7����M�K֟�i�6Ju��P8Z�VHk���>�*��7�k}�٧�����+V��+ڸf��Hz��3z:�~����|�+wa�._����Q�~��p�B�
ퟛ�cz�$�ʮ������k=�*�X�g�ZOD#��ܹ]s�����x�����tuu�G�G<:9����Sl�tlӭ�V��W�p�mM����k�m�r`�Nx�/<swɢ�p��=�����H$FH�ڴy��^B�*)�pX,`�����cU
���۵J>���8ѿ{�����_�={Ù'�+a�q�ɉ����.�2���>��i�����4�l�3���d[���r1(	�HDp8��h���>��3Wä�z��Iv�v�z��ǟ���X�b\!�e����ی���R����"D"�)����#ÓpK��c7�z�ҥ�֬\��h���冏^}�Y��[-�Z��:�O���X���g5=���g�Z(d3F~��*�ˌ��ޯ��uwu~��X�n��K�����o{��������oY��u�Pz�dW�" 3��$�s%���([T'��LM�I��ٱ{ѢE��/����0���o��������-��ϗƧ��]w�͟��7n?�_*gd\���J���~��wɯ�����m��ф5u���>yۍ���J9�_��? S�uv*�㐛�d��|��瞃��$Y���k.�xú��|e4?���!ޞ��E$���t^��k�=w��E���8gÆ��������ӹ��{��ު��>�³���o�7\v�E]�7������^�1�*�E�D݊�_�ˋ0�S����_�-[8~4~��gV,[r����C�]:��7�����h����|����|���v7�ܳ_�z� �O�����º]�x�=��3v���G�*SҊ�hpҘ��3�T}[[�t�{��?����㎫��8�(sZ~@X��;m��"ܿ_�E�]o�ٱcGc��7n<�m΂'��20<=��c�K����J5V��0\��+?�b�Q�"�?ኣ����{P�����̜�l�&K�1M��Lq���E	wj�mfQa�D�G���!�WOL
��+��3��s�£G��i��u�_�a;n�{�����+��5�Y"*���u�7��55596�,��FbLc��1�܂����0p����
�ZB�8<?�~�z���b��q�W��;�Rb�I!*�����7ê��'?�ǒ^&��K@�������uk)e��?55��{�!�h�L���{hm�X��ez�rS$8N��\k+N㎸  Z{ŕ�uwwý��T�3>>X�o�m^�.�d<����%|ݩV�-���xP��?�9^�&sx��K���BƬYZ�Y���lWF�a�y�i$����E��)|�MNg1
}G!�`��#T�moo��G>r�9K{O����	xN�q���/�P�맣T�C&�*%l�<)�5��b��%]Ś����S���/�����~�ߓzm�$e�mI&�+��\*x%^:
bL���
Ņ?�!lϳ�,D���[�W :y��m���2����?���1�Z��=�J�R<�׏e)�,.�����'>��Pޔ���AB�`"������~,�0�請�]>�~�3�N�㝫.��|�����`f���Yc,�)1F��'��E,2��S)&��67��cǎ��џ�|yG���##>b�r)�Z�s��R�1��3~|�v���D2�Rn��Ci��֭���w<�R�tD�Nh�inB"���aE����j�)L�C�Q��uu���~(Y���c ��u���'G��Z����-n��\��ɕц�o�R�1�6��>V[������d���J�, �^}�ᇿ�~XM������Z�\C4�����e�Y�͛��t���}��R膁� %òw� �dHTf\-�������,�ѵv�?�gTG?��8q"�dЫ�5�k�h�)L��,T�Z�|��EKX(���(���d��jTEP~�����K�h*τ��?G�^é�~���P�1�[�-+G�8t������*/(�Ҫ�fXx,1?c����ú2b<�M���\ڒ�H�2%,��V��j�U�OLg��gK��3��_{9T��$>T��UJSi�Kp�t���;W��wd�旱�tͫT�S�QL�D$�ېT"_%��45�3���H]cWG疷�����1����U��\�������_�
k��_���U��i.Z\���%yAR_@𷵷�m�<p�X}�I��GG����[�:��ޗ�-tvt�HU���(d
!�4�V���p`�veq&���m��qybb�v�D*^�K��t]\j���
��P�QRXŒ��bՐk��+�;c�=�3⚷�`]T�
:e��~��Jiޭ�y�1�jP��|)[�
>"�� v���+ˢT��^}9	ݘՖ�d[+�ή���-W�b���l�$�8��LTDk�bC8H�il�׸���i�eX		�UdI�ݚQ�����\�.8[w��?1�'��u0Ӿ@��+=�K� ;�JD�TH�"����6�*am�LN,]��8ŬBKkk�P�g�X�b�rQ&�cx-VɆr�Z���F�,dV�����*�s�㡶�D,��֜���>��O64��#�����hP
�W.]�ӽ�G?���{O`�R�V/�
�+�Xt�`Lp1p~I0��O�T��xA7��`��U4����?r�U.Us��?��V��eQ���,���xY���٩J�,�(I�Ǔ�k��T�����
��m�޹�ҋ�Ι�	���F�����C�efj*�Z�0QC���h�)��_�p�]������=���m�B:�)�T?��`��a%�n��6�ͽ���my�C�Pyf�e�b�1�ˢ��j�+:���G�r���D����q�ٕ�V�z��_|�/�
�V|��/�I|���HcC����4���٩�B��_��W}�&J��'J�5<3;4=�������o��5�\p���a���Ζ��iŗt\����?���PթR������ᑱ�q��W��?z��Jc�q:�����y���V�[���Оg�zzrr��.�����'�hmlB������` l[.�
�%J,��#�M�ƦY�j���	� I��D����7��ֱ�&��G��lM
j���_~����5[�rA&7+0&R��ۢ��*"��h��ۿ�%�"%�hK[��hET�xJ���n�\ޤ�f_�6f��c�\����9�ʽ_��f��cC���J��ߏ�Aɱl��<�w¦,T5��*����"E �u�s,�a��Ȭ�b�D��4��1 D|�0K;�;g�\�K{��z,�Y�)�����Uy�'fff����O�Ta�R���.�������	w	�s�R7~����&#,�1
�V�5���/�h]��+W��m{�#�X��aX6lعc|��:����Kp��C1�5�Ͱb��V��R~�#F-�J!��"@
e��MB�����_���.\X���{%�P��3&J���8����%oG�� �^����--���L�S"ؠ�*�
��«��c�gU����c*�w5/�����hL!:�<w=�e6��c�\���t[@`�WǼ�DX#!$�G��B�"PJ��Y�X�̥�V�n��ě���׭�G)�`Oq�%W544�+�3e:۰xF�R�l�r�PjT=�T5��
�Ѻ,��b��زeK.�}���z��[o��� �v���r�><��NW9xz ��5�R9�����n�l�!>묳,X�g���E�Ur�L!��Ca/@�x�B���|��;��pa�(K+2�q��ę�,�����w�y�/~��`.UŀG��%}S��I��U�ZՍDB:�Z5�;��L@T��OZU�G��(UT+-%�z[���!��t���kvu�%�쬉���O���"�;�Hf�yz.�V����l6���x�oN�Bc�\V)��4w�zxjzӦM�_z�����F$��m\�v���w���UO�U+���)� 2�D�A`1�\p��Ey���?��/��=��ƺzZ�,ŋc1���I�ye(���W���{(��H�	xX|w�撢D)�Y"�P��f�P��+y�8�O�(3�[E��ğ\V�e��W3�it�H5�	:�:rx��_F��U�z�BRD�hU�Mo���@'$��$�Y��{�����������֑����x��+�R�H�Xd�m�6L��8Q���	p<���!~8��C�`LԐ�W쑑!���B�
t�t+A���CrD�I���k�YT+����̂�s?�tv����O��	Z`�6�a
����d��.	J�p):z�E��im}��	C3�+�,^¿DC��"��TC��>�J�n��/�)h��� D�e�6��	(���;�)�ѳ�l�,�EK�e���njl���BW"^wbh����ZZO��海�3���Q<�dzv��s��VcSJU�|%O���[���W{k��E�T�ϧ'5-�\vI@�2S���$�e�V�M)��C���4]̐���DR�k�H@Pe����≘$��V���73;��J��&����I��R����a,��T|�15ʌ2�#Iq�W� �e&%
ׅ�Gk#0�����Xzb����(�7�n��{��J��f�d�|2��*���m�&$3b��Lz&S6jr t�x?����7���8޷z��H(�����پ��;S���ҳE�����z�ƫ�WT��d�4���GScQ5 �	��Y*d���eKS%s1���STu\5*#��^[+�<�UmQA�Zb�<���� �k���K9��*���Lϼy��W]~�蘪�+�r!�E����?�����N(�s�LCij
��1�."�N�`ȇP��f��j-�-�b�j՜����1z���߾�����cw�q��Us-*a����jX��JJ����T��f��"(��i%#��.[��
�x�U�/^~��_��)���k~�u� ��T	�!Ѵ�P �e����A�'����jn���^�IOs����2><�ȯ~}�]w-]I�e��K3�|���Q���d
�ZD_�bp��U�	&�{�!�h�;��+��Y�,��$Ebg�Ys���z꩟��/)=�%u�9�\�����?�؟^���`SG�c�N:��8ǧ�}���6 �H ���?�w�����Ȝ9-�T�j��J�+.[���L�v8��Ow�U�9L��*�Z���^��B�X����#�Cqädм�544
�᷸B�v�)��XoU;�j�g&�.=�k���h[��#p���=���E&.�jh���e*�r���`�U UK�Ng��ʹY8���cp�*oG�V���C��+e��X����*�G(�З�nl��T�̛7��1��^���5�QUg ��`���M�~U�Ug�B����Re��UV�e_�&K��5ic?07��:g���SSyxH L���)Ҁ婼 }��������*���T0���5��m����v��Ղ��(��	�����X� n0�,!2Ly�&�-xB`�T�,o��9����kȏV!���]z��x���=&�{n��<��e���]w��w���qL#�tL�/�u�Ȕ���@D���+�@�kr�9碅����X$��4��]�e��ds��%y�|N�u��j��0���9&�'�馛�	�E[�I5(�G��o~��)�� W�o��d���à d.�t%�D+H����L���cN�۝{J ��e=SS�۷o��[��A���w�}�K�""rb�	0@�����m��
�Z+R�d��t����Ȇ�"^����)��u���x^�&�X:+�c��g�CәվL]v�e�c�:��=
��_��x�1�t�
6�!A�������szQx�ux�e˖����n��t��M�����^��ε*�-��E����v�&�t�O�l=Put�ձ����^�Gc���k�A�����@<7�|���������0>��MM N@���,_��%P�j�4K�R������J�Cc�=��u����T.ǽ���㓔p���/��bcc����9��P�$1T;00p�豍�~�K_z���ҩ�DBx(����}%�T��Ÿ_~�y�{�*�S�x�g�74y!���q����d�F���Q����]{�5#ǩ�qݺ���o���?�5�,�b��^"<3���<� ��=�'a.�###�v���n�{������������?� �����|���J�ܳ  ���.]���������+cybL�T���Lf���:�Be��ޡA̚�U�������,���7ޚJ� ��:����m�J�J�[�{��m3�Va����<���S��fyvs���a�&�d{�iˮJ�����/F��8�F�l�}���e�<�][��r)��[S�2���	�iٜA\�*�
�eSwm�8A�L��(��(x��"�:�l1 kt�R�j-��)-�����,��Ѐ0;�m���{�w9�d0T���CB��3�[�|	�Ҝ�_��ے�O��O=�s�΀��o��3����EVl����SMR�c�N���M�F,9��2��UL5���)1�v���b�r��N�$��w��X���n���!8���|��c�,����tU�h���Q��\�l�y�^�x�9�Tb����q!诒t[�X2'�6q���@c�@�9�
I��O*����w�=49����gy qUk�9���}�-�y++�]�MES��FPv��f)�_�i��2��-�-r0�P�MN�⹂�u���߽�v�m=0ps����}%� ��ۻO��b	Q@�J`0ކU�H%PL�(���yEU�z	���Ɲ�ߦ*\�������w��΁�i}���^�y�c�U�e�Y�M�Zq�F�r��)d�\��gh9��!�#�sLi��lY3�]�e\4��M���^%�ҼH��n�/ʜ�r}S�����DB�O	��Z1��q�B��B���V]E�B���>�Z�삫��x��en��=�F2U�qN�������ȢE��n���y��EJ���R�*V��0	��NKkS4���w��4)��ϕ+���솳|l���>ۅ��r����-�'[v�+��jL�T,K�ٖ�M}�˅%���u�L���ʫW�p5֣��3��������L��+��/�.������U�޾}�)�H4���=<=^Ѫ�h�9丙BE�$+�K٪��M	n΢%?}xC��o9Y��ӟ���n��l�d����X��K�=������&��ё�ŀ(Z���K��u��p�u�W<8���LL��i�f�#�ّ)qy59U���K��/[��\��)��`���D�v͍7^K�TDflָg7���)sRxx�d�܄+W_ݓ���7ܰ������o8�ӓ��7��l�y�DxݺyǏO��w*��/rEUI�OJQ�'���H
B�b"�/�'ئ�&���{{_޲��k�=�˱��?���$��?�����zO.[�z��{���O<�ĉ�²u�����I�̍���[��f��͙J!H�5)��I^	�1FAN�S!�ɻ��wG���;m;�Wl�o�߱�'|ۭ�N?�K����S�<�X[�l�p@M8��V9
�+�0۵`X����&��P6 q�%�A�f�o|�i�$� q��;���K/�|q�d��Xi��kB�b�=��O3r�4/Yi�s�ɝgt7�J�y2���="�C�sr,/±O	�z� ���;�P0�������=P���ޢ�Ҁ�T��Oԓ]�
�O\��r;�'N͉�	��0��^���klj8.����c�
��1�{U�ރxE��^Q�6�ep�"q�n�Y�ѣ։�A�s� �E�T]�g���L`Bv� �T��w�y�Y��������,��(�^͉0@I/�y�F���xdtT?6p�v��!�#�v��eh��Ç��كA�%X&����O���F�	"�p����33>�HU�m��ٵ}���6>����T��������_��)ց�HL��g#<�tb��˄ӕ&V�J���h��?8��3�d�ʂ���v�<A�`��y�(��;7�������6�d{ct �9/��ʹ������G���G���Y�v%V�X�0��X�d��ƙ�!gT*,RF���Y*���e���%Ke�)Z�x����>@�^x��ᮍ7���wh�=�� ��ըN%&���lס��@��Gg(F��ʓx�$�hzroU�6 a7w��r)#�+Z�J�� ڋK�<#�̙\}��j�T�&=��dWx��7�"�΃�����@O<��[����Q�z���J��K&F�Cwg���*r��#��x���#�3��s �@?$��~5ຊ�<�$:X�O"@��k�����S����sd��ݲ���>�Y����l*>y�}�!��s�r��(�Y�⢇����l�222�U���q�bfv6�Ie� >�x~'��?�)b��.�x�e++U�С�W^yi�޽B0�m�㾅B�SQF#�D�P�P���E�A�bpp�9^�����r����O!����+�d����~��_>�����o~�{����F�{㍷_{�d2�99:8� �Ϫ����`�NOsC��cx8��/|��5��W|��;;;�n݊9y��7���3Ϥ�Fj��Ȍ��8�IMW��$�[��g���:soa�kD�)��h�y�w����"эp^R����[.W#�.�����Y��Y;ͮuBN���чbj�T������D�L%
x��ʖ�g�<�8et)D�Q0Y$�+)��!U	����HcfpFm��C��<L�S,��%e,1[@���W����-I�d����o���^ܼ�U��$%����wA3^}s��"���@��~u�֣'N�K���	��
����}�ڵ�h �U��N���dC�08����Fß��7ˬE�u>%�	���/���{M�Ĵ���#�����̲ͱ�Œ_l^:9U{~������Dw���\����'a�w8�g>�df�<g[��餓,Q_P���0��J	�����)��r"{�b�B�+�>xrώ��ׯ�xrl���Z$�e��n����xxDb���frS�'��q�)��^y|���U�B4)��̦���4'�'���\x_$�����cci�$6]cl|��(sh�o�X�C'��{��I�T���s��<Id���b"W��t��'�4v�)�xk���'��>"�H��5�|��(H[�c�_��,F0O���������{������S�a_�J��5���M	|K�Gh˵lͰ���+߰m��M�Z��*�;�.!���}RU/�������N�-�@��7Tkm~�a)�.�~��B������O(�mF)W"g���-��b�p��w�a��"N��ֶ�h���@MB���.Eg��� [�p��=�³�n�q��Z>Kh�%qu�����36��dm64S�;B(ـ)Et�#����G��L��V�nذ�Z"�vB	Xr�q���b�`����l��}��o�b���g�?���oy��B�$h\���4��ʮCG�~b\���E���x�{����3���i�}~�_�} ;[�U0���Y���s|*��_<2����r�!^s�X<96�����
?��A����hKK��#��Ͽ�iӋ|!C�{?�c��`�^{�����X4qbpdplb�k�lhj�k�H��G��*��`}>���R�8����0<����-����/��'R�X�s����g�96�>�*(�z�x��w��d�[4[�C��ʚ����N�9���BI3L@�`>W~��}�"�^�X�����f�e��e^����k���5��g���{�����K��0����'lr�9��N�xi6�8H���*��Y!�� 8���J�K�E���<��&�[��X�Hù�. nD�j2�.�����>�ei�b��HI����9؃��j@m��2dp;��-,�l?�E���jթ�$K8J�`V	g!j��=~JL�⬆�$�$`m�� �D�WvK�#.���c������8m�\o�d��a<��:Xf��f�ɖpP%�Dqw�څ�)�%��d3m"�u��eۗ���,�D+1���EG�3�l۶-��z`��: ��kH�� $����v�UF�ĉ�w�)KǢ�)�%O�	O�m�28�|�oa�r��
=&��^2>�����]Ԍ�φƠ� �j[;U�64x���.IpY5A$��",����q�"aI���#�Q��^^�yO��mok�>��x�ma��(����IHDXj�T����Y:�q��#!'�FE�c��7oEp,;��VJeO����$:�@�Wp��}tJT�N����F���7U!�d"��:68������e�jJ��
<[e���x«�����C�z����AU?�B�t��mz���Q�R!O� �ZdY��+~�PA��"��SӀ��LI�;���!��Ø{�"�͘��5�S��e�֘΄�ڬ��QF�\;�Z%�ϑ��N	K�p����'l��=�ɖ?1���Rֹ KC�,ç���8�+7%� ���^hK�%J�`�Q��%�Y��CL�E�o�γ*����V~C�U��w']DBv&����_y������o����9r�ٴ0�.��h֣G^�H{�z��"�p�N�["�r"�A@�.��d�*�fCI �S�tr�к~�����}�c���Bt�  qy�ȶ(��K��O��~��%�1FKb)�K<��'dAО���j6�"��!�#:���� �� U��	l�G�Z�jy���PP,�i�U��M�����h�h.+k*̔|����$�5ͭq�T�O��Q����u�.Hl�N�bb^�@��0��Ua�I�Z��Z-�N��r��#�J�»��Z���ߨ���lADe^�U��Aѡ(�d]��N�N���B ���"�3W)��Ĩ|"��T]N�)8U�w,E�e������l_<֬���_8Fhc���!��{M	���\�w�������d2���8�����H���2�)��h� [:6'��5K���.bp���Q~�V��,;J豨���"m�4� 9������MW���l}C#kI ^_(��b\:z����/觍5���A�ozz@�I�=_�]�H��;q��c�jqʹz�O�"9K�O,��	����q�dz���{(=��2�i^�L���A!���NG=�o|�*7::k��|a�ܹ�i;�_��
�أ�CJN�5x_ô�T)_�"����4eb�-%�b:vd:z�*a1 c���	]"/��j~����t�Qdc�P�pJ(ԡ�F�FD������W�.��65��CuXU$�,����ov�T5M/�fgn�O�ef"��AWd�	Ūv�r.�9��Iu�*���������v�)��X�>�� �����hiF8��N����b��)3����׵�33V�*�+�JEM�L}j&ah&��d�,��ɖ�˼��W2�H�1G'�*�Fu��(���M���ۖ�s`H���e��LY0�U]��AG���+����j������+��,��@rq{3��-�45�)J���|���kZ.�x"�667�f3�BYF����br��ã�g�.�$Jg�h�5n,N��,�-��Y�b��[C)�S>�)5��S3��&���LM���@5��r�B�#Rj>%�ܜ�Y�����E5�
4�����0�!/�fC��
0M�'V,���=��}O�����w/2�o9�����y�(���{���[�L	O{ދB
��hU�q�A���J�h�B'�eA�aI��u�F1W��ܩ#
F^�
���]����O����+��	� �.�
��װ��4��!��d�n�N`4,Ր?��egf,��I,�ёq*�e��^Ԓ���&"h�T�5���V>L���xL��)1�L|�N�xO'P¾�JKSR�Q T��c܋r�|�7\ps���(���ۄ�_)��%�a����dX�����G���
$cb{\���VT���Qλ�yE���(K�� �OO�c(�N��N�4�$�^�����|�&hÄI�x���˃�z&����@�M�G�*H�R�R�V�%̇��}����غIk;g�y��P���?�H��-b���R��9��'	1�P�(�������So�yGA$��"�^�*�Ɠi^�h�"�+�yJ�Y�z�UjԘ�R�]��<?�Aا��>����7�9���Dk*���~E����*�W��x�JO0 hs>_�xUѫ^��t,�UP���@�"y��y���^E�Ǥ��c�Ä2-ū��?����}��)%a�bu������]�Pf�4�0�џ�����h��� ?a�f}S:
_�T�h޲�<"��CP*�a@o������h�#����kL����^-4��m�+0Zcj�Y.��NY�r��ug̛7��SM/�Ϋ�Ã��d�D�4J/6t�!
��n�GűT2�N�L���2y%���h�_f�T��N=�&�����뮠�塉����%��3C��i%��'�,��H���ٻA6+\Ɓ�R(�hY2;}�ج�1�b"��ƭuS?���?6��Z�����&ڰ���L�Q����O�@ݱ$�ᥒ]��g[���i��$�2��]��wYވ�bg���e�.��8�yK}t_V Pe�6�V8&)#9u�����;�vʹ#q"A�=F�]��P� �R:�7L��dR9) _n&���.�y�L�j�I�©�-�Ґ��L��4�jLRܓY�sKr`x���-�jj�cY�O���%�P���T�����Щ�$Y߀in�X�����[�\B_�~��5�`%�ߴ�����(�F��x0�� x�.[�^<DFST<{A��>
��w��P��d����������R�X����=n�ȥ0�'���4<��Lz�`N��tŪS���x��CdtXA�aن�#~�݌h�𻙟N������O����{ѹG���W��8q�C ���$A�̂�$�J�S���J"�V̙�&�L%C��F�3SҌ
F&��i!�xb����4j���
��cW\p�@p��:%R+LH	yҹ�V\����כ���3�4�?���{��904Gw����8w�|ڥ�J {~���s֯B����K"�bY:��ǉ*���}��Gݶ���=������eӴ8^�� T��9'Z6'Ҷ��l�8�7���0 `�HH��u�V���9��dԒ��fVk=04JH��K6;~7ɂ�2��K�&)����K��]�J���J�$�E�뮪����.�\���=���VYJ.��U�g֒hl�j�U����G"3�U~��f\B}s���x RgՈ4��;d?��Jj�\c��@A�f�m蕠꫔K������:�
%"��|�t<�/�9�Ĉ��4qYr�ZY��������`l��Ūʵ4�4��t�UYE��U:�Bw�^M4)���pd�U�D�*�f��o��ꫯ��u�P8ø]]�@W�<A�H((�J�#��P@���ƵK|���tf^S]w���{n4��j�����m5FU�� %bTL�*B��+�D��Ҩ>?R_����)��u�1,��P1��Ym�����Cd|,�ģ�`��
�w�9��C�Ng&���ato�3�I��O1��S�?�����h�mD�J�'(a�_�%j���{�L���S���U"eUپ�^j�Xlg��ე�îL��n���w�=eK^&�SN��c�A����xt�^�+��xI��H^VC)�!�����}��_��@��ގ��z5~�÷�S�R���0)qǤ�:���Z���t�
���\T���*��'�HU�x**/�{�9�y�~��-x/}^�&�=e/p�P-��	PE��O̲B����*��\��}�5�,]���[o���k�3��F��ƘS��/�O�M\�t�ڳ��:�S6�
z@�
2f���B/�V�_��c��U�Ĳ	�J�bĩ��a�x
��Zz��$��A�R�e2J,�@!ha�X�#8����^�ҍ�ݱc-0��`c��@�萫��f����?���B!�UW4��
�-�ܲw/;�/��]c"�ol����R�.]�n,��ݹs�! ���S8����QHBU���f!? qv�w�B�@5<�)�QF��]9;DGy%�EBB��Cct�088���	�O�8���>���(PkaJq��vD���)�Iůx	u^1*eı�[&,E�NJ�R�5;�+�PT�;�D��p���%�}\��Hi���V��/�be�J��UϞ::f�u&���M/��-.�	�����ӌ#"&��d�� �����%" ��).,P�G�Ȃǵ�����b	_�d�x��HL>�\�)= �aJ��ko%�Y�	���x/�ܗ�̪�MU�R���vb1��]��v�Ӟ���i���pδ��،mml60 �
Ђ%�U*�T�*՚��{������#"�J��ۄt�deF�x����w��U��/�^������~�믏d��N���d�OJ�����-Y�h2�馛��O>q��B��N���355�_>�W� �ȃ�b\�&nض�@\��5Q�B�`Y������F�`�۷o�������c��]zC����"�q�!�?��1.��oG�Y��A��fT9r�Y�`�H�e�XҥZň�l�^w��2�T�g0��G�1�oZ�d	wXY׭ƚ���f����S5�ː�!�O.��F�;qh@"���:H�R���cW�4:,�)D�aX�2#�����P����冇!���(=���T3,d�Wh�TF�s#�d3��Gd���~(�f$aJ+aAZ�z��ӥ�f��9"?d��������h�Ht5 �r�P���@хYrlx�P��(��� ������,���t���-�)(�2�TM��1�,
m�vE�8�p��!�F��'�k��n��Y[�dZ�2y���-�=o}h`2k���w���1kb��?�w)�}�*?=��f���㨜���k/E�F�)a8�V=E��8�"�w�g�<�g��W\n[�={��ON^~�ջ���F�Tl5�4_���e����">J6j̝�F��KJ����Z
T�	lT�!�<��qr��-w��XY\�	�G���v|�}�4��	;'$��?|�{hs~����p��#p!����r�-��/G;M��>u���~011��_	�)���혚|��o;�:t(�FzԔ�j>7@�l�Ȼͬ�r���Q�DOZ��Y5h�4E��*���ڹ|&����Hv<�FZrei);8�����,I�z��`HP1u���
<��nj>v��z�o:ER����]�\�B&��^�@�`�JYp���ӱ����'���0Og
��N(�LL�-)��W�/>-P�������0�� ����9Sá�2�L��rp9D�:�q�TCZ�ܨ�^%]1tS�e�P0��P�4 h��t.$v5�U\�i��Xt�DV���	TXj��]�~K���<v������;��WR;C�SF���FR�,�N*�1�T.Пx^�;���	^�̏R/�c.���O�yZK�����g	��y�Ɲo�[��ִY+�A+����*��_+��I&��_���lC�RKͲr��!�)I�h=���fK�y�`+�oy�M������ˋ^I�l[Z�l��sssG.�B�23\T��"sN^y��/�Ԭ�t4A�A8�XI1ovjk	��
�0lxX�B�Q<Q�r���.���\�����BO�ɡ�����UR�+�N��܃��H�5K����E�"B��4��JR����i�����xѩ��Ԯ�:���l�a(�A�Ȃ��OGē��ku�S�b��͘c�°`Y��Ò�QV����?�<��Uo��mZ�䮚��Ν;�+M2Z�eP�LNOヘލ<fX�������Ǉ1/W��sr#�����;�0}#�R����V��O])�I	te�G�E�L�Z��C8E��מ��q^]A���6���2a���wp�[l��2��a�<O� -�95�B�ܓ,jW���Ȱ5<��D+�ʚ��@Wk6A���8��B1G�=��2rt��f��R0�H�F�n��&9��]W,�h �
*�{���?�/�5�徱�$���I,X}�o�vDK�Du��[�inu����<2>���C���Ze�� ȗ2@yL�Y{���^�^�N����I�X�M	gy빱Myn�P{��G�C>G<B��|��-�i¥��Z\�^k4�kC��������R|CH���:�R��w��=����7�yxj��<�,�*⥑�:@�~�!]my�#�HŇ����J̔�����dD&�xtt͔��������/��.RnM1�ں��W�w��~�������`��M��Y�v�<݆�2K����Ӎ=����ǋ�[+�_�OOO[c��OuÄ��M�أ_��o�x��ݨ�{��r�%G��{��f�޽���+�YXXx���G��X9�Y.K%c�6tvrB��T*���).W[pXȊ'�<���d�g�\6�"�r��-/R�hlY|A^Ai��`%��ѤhI�ac�-\_�rj�?�E�"'=*on@��a�%6��zs���R�x��8����(��1�Ng��(#pKNF©6tM+��~c� ��sH��U�?�PM���U	h�s�U��u��}��ٰM#|-i�qc ��cs}!�����]�����o��\_�y�{�M#x�#O>~�8<��\ܶmbv�<Z�FGY�8�gٮ��ܒ*eggg�=����͛������][�{�?}���g���%or�Y[��)�/6X�:Pl���J�IX�)̜#�9/@[�UM�Y1N(`�3$��6U/%h}�����֨2�^�]yńx���ת��>����CG���aH��WD�řo��m���`(0l��&)�|�+ 1N�-�nwyy��s��ܳ��<[[[��͊�m�$i���Bޯ��jI�S�h�Q+E(=�m"�+V�l)�/��}#cy-7l��l1Wtؑ'=�Р�>2T�'�C�1��Ӧ��,�}qz��փ���� }S0����D��31�����r��O��	�X��� ���	��k�Dߟ�y����u�lʱ0 q�m����&������q +����t[j�kA^���t"��u2�Kh�lE�٦(!I�yJeK'�a����EJ�?~�����7o�6�.���+�ȣ��\����~�ُ�[XLKS���q�=����M"��uSJC������x�mJ������c��c��Z\�h)��%0%�����n�o~�5��e/\85���:�R��Z]�h���겖�vn�?��O���_8z�h��?�kWNeVv���1z#F�&�-�#�^�7����ښn�J�KC�r�)�����S�uB���-`"�A�ozӛ���j�.�O\/���6Sߵ\T�Z<��!,����lٲ��pD��/�խB��!W� �Nw��q����������A�d$|#��:0�ߌ��.4:.��+�C����<]�<�<X\�c�+mPԩ["��G�qC1;��D�q`���U6H!�6u&Bva�Ϻ��n�Jh��v��}���'N�����@BМ���s ��<3����ٳ$��vm#D,Jԯ��
�ۙ���SN�bD���}HdeQ�1��A��6�yn�b��-���DļO����J�n�ȐroV+�O��|
U�bH�`x��C���Y}0EN���&��~��-�xv9ϤEii��y]Fz<����Nf#L��T(�Yu�*UR�U.��b奎��C���+bG]y�:LU_d�&	ǋ̪�%�U.�y^���c/*"��vlڱˤ�$�o���aff��bjjJ`�nAȊ�xhH����P,TڙI����Cq����ݳ֋0bi�'d��/R�]I�����}$��Z#�f"s@����=��)�0���t��G �4�}*2�PRI�B�ǆ�;��A0��Bc�v��}$�Y\������珟��D-Zj���Ԙ6�<#D�!صk���Ѫ��5����RB�.���*Ϡ��߸���s��!*����k�E.��Br��x�ȑ;vl��h{�f��B��1_�����3��\ja��g�;%�j;P[l�.E��R8Z�/��K�d������!Z��ju���[�t�@B��I1���z�NL�5�V����M���&ZK4�_����c6�%ꊎH�ʛw(Im`���`���R�:�X�*&s�?d������8����͆&6�_1�I9|�,UD'1�4@�l&��h:���ɽE�"�A*>9�%����N�_��L�T	��)���HA���n�I���ά��eH>�#viS�����JNW^��^��W�6V� �{����?�<�D�?{a���?~�?��تKǞ�IV�o����z�DPQ�s�{�͙˫+�����U�2	 ���_�x)��??���o���o�GJ��I�OONl��ٷo�m�����K_>y�dCɐ1(����Ωݐ��p��c�G%�F�n[�&4"j'�.<��z_�rruwN�Te��^ ���{pH29�9n�.G�x��9tE0�]��I*tY,��9�:!���#�����2j�8s�Z-o����1�$�<N�D�XVtE5HS�P����h��i���!��U{Df�nҭ4m���jn����X�H�`���ܚB�s�AGf#��C�56꺪��%PY]U���=>��Vب7�J�b��{�{�'Im+w�<��'
C�V�uQ 35��
O��Q��e�7�'�*d.��h#��f��r}/;:�k&�	�F���6�p+$5�3r�&�m�/i�pIv��b�!�����~�
LkHu�o��ٹ����������s$q��S������?�9�06}9AǤυ��Ld��ꪎ���/�9t���q�?��ĭJ\�X+V+U7�r���d�u)P�xm���o�a=������9+�\�Lƨi6"��r9L�򕯜)~�����ɡRq��+IW=�]���ڮm�f<?3K�?=Z�܍U��~~W��P��/��DR`�;��<�jzz�P(
 I���z��L�$����ٳg��[�=w��Y��:��M�_���Ax�3XX����_��j��څ,��!��+�u�B=1zqT ���������ԯ���9P�{�]s˾���)Zp�"-�����w����3�0�O$�6��I����|��n;��쮽���o���[���dj��wߝh���O��]���n^�o����,�_��[�:��{���[o%�>T�K�B؄ ����_��n�y_+�uM�����,��5�ΤQJ�h���� 8��8B\x#
�<�z�Y��w�� �@��]��H:�H�rw4<��Ax	K�+��L.��22�rij�o�F�w��n�|+d]����������>e�V�L:�%��(�Dx��"!��E霨F�+ONN����9��u�?!�.̗�O��Srw�*��L8l�޽��3�G�T�#Ae��N�#��-��X���R��O�,!{ݬC�=ǡ��M�/�w��m�h9K�J�3ƹX[G�Z�Mڻ���U�7��Up�f�/)*ٌu��%'E�o��Δa���P������ok^}�{�C��u.鯪��'>�	RS���u`�΂ �'X
����i��g�\}��t�\d��:�Ej�0G�_\��c��O�x/����=�f��;���w��]�����`7Dp�n�����+�@'�$'�cE�S��tT�j��6�7��M��ѕj
CSI��7ei��0�璭Ξ>6/�_&#Ky�����|N�+�5Z^������+�L���WW֫�P�k���!j���?�)a��łHl������1��'H%dE���� ��(Nخ���Ic)B�=�B ����n���C(��B����Z^)d�k$ ~/EL,� �:�)�.f􊩷��}��'�E��VB��D��t��s�+���j�hRm� l�ye�诡�#�ހ�
��N"�kF��%���'�gg�Z���2挓 ���t���c+߸���<)ES��w��J"Iw���9���߲�v X��hy�����_�?�,��w�7��Ç3����3���'(�5Zͺc/,�4OO`�Tum�U��W�)���Z1�	��l�9�zqJ�]D���d�I!���|M&��#,I5�S-[�2�:�e�&U%��;VPq�e�i{��l��-L�FS�]_R5G�=?�HUb�)S�,MM5���O�T�����$��ɶɒ�װ�H�äpD3�~$��lfK�W �!v����;+��VN4d�K��(�vnd��8^���q0Y�ހ��<�@�(I��n9��8�@�.	eH>]�����2�Ra..�l�:M"I&��2��$Wuf�.�����?��Hd;�P�]�G?�#q�PG&gT���v�7Ӂ�i��Pp����e�rDh4�r��֗���a���,��ת��Ia���&� ��S���ڎ�� �b�r��g�'�薙�ڍA4F�ܴ__�gx[�l>t��ԑ7�p�տ���|�?=�|vp����֠p�u�v�T�KJ�����0{��n���>��*������������gU�$�1kfQ��$/��F����w���~����P��W�1|t��ب���K�����w�����N��S���JXsK�m�.۽�رc����Z���ZRH����5]ܢ8���@�d���º�Gi����651A�ޅE�B�<�Q{{niI��[�Wj!�Cb�����T��{Ҽ�IvY��u^zM񽈢v�x.�Ñ.&2��v��� ���&b8�x$�]2�@"���{��8@)[.W�7��D䗖跭���gO�ڇ~��P��sR@慅�W��5{���F���ɳW\qſ����vYxl��p�(���7��ȋ��� 8������_8z�[SSS�j~a��]w�566v�ԩ믿����k.�NLL\h�ܕ�T�]�&�bb�a+����P0��� ;\��/�:�(<?��F�� �f�=q℡���JVJxfV��	8�B���4�p ��P�A�B2/d�ě�D��E�]�,zh{C%b���E.��|��tvRL��l���AT��dUAWG�
qR�<ql�֙���ZY�c��r�\*`Py��*3S���*ǽ�$w�v���CURǋ�c3)��E'��)1H{�E���A������m>0YT��m,.B?�\�oOOO��*�Ϝ���&Sim�-L�wS��6�")a3���!,fYH�.�SK�k5�Dom���?�����뽧����?��'Σɋ]�<�$(�8�`ɜ��ɯ]UQ�p��NG�梳��z}T���Oo�+��y�.��c��=g'���^u�U��{��݌�=�V�OG�4�b>G>�QT�P^�-�v�N��B��C���������/	8H�0�mI��*P��H���ǒ�zRLb�s�cǟ D5<���
=��r~�L���$gۦ�90���1�V�Qo�l�̉'S)7���*-o���؏T�ǚ�A8"6�1�F=�旐S"ܺ]���P	@6H|���&��
�
ac)<�<Q�xĈ���Q�@$�N��'+j{H��`fC�$���I���Ȋ	��xk���S��"���ꑙ��&u���Q�D�,���5��3�$�%�J����W4�,S�B]Q�ZP�뭠Ī�{�$w��\}�R
ы�t'J�D�Ac�w墡���������Ⱦ�C�J��'����?�iy�C�be��Ֆ24��R�ʪ�s�$��~�mw�}7�К�V@�!Vٝ(���[�8��+��~����Yr��8h��Յm۶��o޳s��@)g?~�\�"g���d�څ�CY��R���܈As�_B�W�bE��#���Y'�$QS=u��+Y����x����!�k��V��o��VZ#�t�[-4Ӓٱc�4uZ�G}��,����*9WQ����RPv��7C͐�ֈ�j"Ճ(��j��i�+�?)�Z�&f!���Ē�PBH=�*rW��z@�`{����@�?�M5�T���,_oxq�o���rN�>=�W��֪k�� �,�3K��c�cc
Xr��	��c���竍E:�k x�����2�k%�꘤EW�0jm�2��H�3U��� Z@��帹F��B�^#�����1����l[���L'Kx4��|�tD�2�%n@(Ec����>NM!��������|�����V�4�j��m4��
�5TN�)b`	Z�`���X*���!5Z��/v8y�����#���������?�@4s��O�h���45O~�/���j���}^�~�}�򓓆�3�2�Ӄ��!	<:?� ,cJ`�W)2~$�_E^L!�)���Ƽ~*J�s}[f�V�d�U����H��8C���mT���*k�n����T'�F�r\�}�LD�X�K���Z����5qzH�H�
bKA
O�ǎ���o&�077' X_ UK�&A�����)x�7c� D�wzܱ�ft�ǆ�ݺc���\�&�/6u=1��ݗ ���Cn#JE'�H�0�H���$"�����^�Ai3]Ki��=�g�{P��[�p_1���٘N|~]����dQF��y�OL7s�����V� :&�K���w�}׮]i⏏���.�q����g��E���>w�Dt�k_�A�8���������������G>�{���p���_��#�<211��[�"@�$����>�,�������[�={vdx�>��<]�����g4�.��j��ez�o ��r��P�`����ѣ�]v��W����z�O��\���m�VT��}���k���h��Y	�ig���7Kȶ��bX��䊹���t#R�>�vIxu�
��St����Ο��K�~2�*�3�޳�C��zp�'?���Ҫ�T<�%�X\��2�G�l��_��'?����x�@XG�.Y@��F�Z�k���HKн���<�)�7;M�n׷�.��Ξ��iA�;M]����	�|ţ1o�Y!��$��ٗe��@�BW�gP�V7��]Ľ�ig�\F|�\F��vjm~��y��L�p?fx�M���m��l�@�v *�)�������i5
Μ9cFh����H�q��GT��}�r��F�
�QT��Ψ�)�K͌&vIJI�K�>��z���i����=��ї����������@@'b�I�Е㝿Bwrau�'Q0H\k�]����z?�t��L��`߰�X����d3�dC#��Qk���6�d���-[0ڍg����8��
oT�t
Ӓ����U�"�/��U (=���a�2R�4���R=8�QR�=K����T���HL���~�S�s�"�Ï���tn�t�{,�&䢽�]^63�����C����$�DS�y�$�bDxc5�ڐ���$�jY|�1:�@���ٙs�Bf�޽��}��뮻n���Q'qw���@�{��N�������kk+k���s��ۋ!p���ލ��~�x�������塇"�`��σ���0W$v?���>�����y$\^�Gf�V��n ����f���/'���9�N����0c�;HBn���s���Wg^8v��~����Qw�d
�L&XjȢ��bA��4]]/�K���j��N����kn$Zli���V�j4
�q�٨W��ֈ�ٜi��^�X e��\t�+H9jh�ma�O�/� ���ѹc9�j��;�Q!c�q��t��7=+>J�j(��i)�&��VS�T�(�啅�>3��ڽs{.W 'h���+�
}�k^C���Rn���B5�9'g��F#��Uo��PA��f���A�aK�/p�)�7jg O$j���F8�2o
3��/e�ΰ��@��ٟ�xS���G��'!l=g{i�r]=AVP%�_�k�N~�jj�f\s��zu�\�v�F���=nlYU��0�;�T���D;��j,��Gu�J�`j'[�ZM*�F���3�:l`�ǜ�D�?
UCW����o�H-Z���e��5%S�.�#��!C��%m����t���*Z��%��*��:�����g$߬�lݔ�e������<p����B���R�&�bm4�V�Z��Jf�ja�	����%:Ƭ��t9(�T��A�9z��B��� �gjj����d�^���8p����ӧ�����:v_4^+�Ual�����3��:�.�UE�1v��Ӵ�'�͝n�e���>;�3�&���u�[	IV���O�Ѭ��������zP?W3�&G����&�ҭ,\�bR�>�-2c\��G�˷-���'���o���m3;�?~��sς%��W�Ս/~�Q��8t�)��m��F���o~�v�V��O���~�p%�"R��,�(ug���)��O�t�MB`d��'����{�����G?�0!�{����?i1�!�%������gN�g����ݶm���~�g�gd�Hl���Y�Dһe��2�ؠ|��Xt?�,�y�u��C�{w	$��+2|V&��������H�&⧕��5Y����^Wke�Dv��,"]���B�v1	Vt!��u�Ś/v��6���9�6Sϲ1�����?$�(;}�=�'1o5�܃:{�&�Y��莦ǧ�c��-ɁR���V���Io���k����%@h'YE���a���:Et���c-_�y1�ƣq��@Gi7ڃ�+�˪~���XAL�/�(�쉴�����8=!Z�UPD0-
`��]��a�࿘9���͔[��	Œ��+�ɀ��B<<4pR���������-Y�Om�� <���ƪ�f��+�W���q�J��uvja����Co�����Zfgg|�:J_�җ�U��F��ʎ�7tvH�*��?��r��y��d>��\��^�n�����M�Av��O �}�?]�5	��3�j�r{ +Y�9���g���Gt�p��f�n�>��є�Y�Ĩ�#N�qI�}��lQ��F�>��q�rV@KE�S_�)�O�v/m7UI�w-�%^X'�/uE��6!L��[���W�4Nծ��Z(������Rp���%p�h��HR�vu���!GM�4�R�������Df{�ȩ	�Y�-��f�I�$X��W����#v��ϻ�y��s�>I��c���p���=�7��uR��+kW\q��7�L��W^���}��f�Z�f1쐼:R�L�&J�*�*F�c�󦮇��פ����_�1ؿ���ɟ�r�׼��U��}���|�ۤ}Zn3ggϝ;Y�:��NhIx����w����0��O��W�1<F.B_n0t���H��	�[i�Ӵ�p�B�H���LlϏ�o�O�1���}�~�i� �^^^���G¶U;7;C6��4�(�n�E
Uo���.m>�L�b��`����U�A��v����L_.�w����cD���������(A����Q��PI��m%��14�\ٔ�%�Y��ld�f �fX�<����頭���Ch:�R��A�|����Ħ%���A�>88���7��U A�I� C�:���HCR�8�%��F�I"�
���NX���u� w�����G�l�8֤T�T͘��{5/"(��UE%�6h4����|�8Џ���S/ZΆ��f����6�U.Q�2w̐��	¾�
(꼠^.����HA� ����/���ƞ�Yc#�f�������e��J���R]�!$i�JCC�gϮlԂlq|��n�jn�������y	ԯq�;l��e�"yN�-m۵�+_��?�GW^}��?��\��W^9�}:j�oftt8c%�>L���FP�?��Z���,���& ��W|~�+���a�t'��&��!�"�%\-S��z/q'0������hCጙʵ��7�;	7����ya���`5ՈA�ڋ���m�f �wuo�|���߈�c���ޯ�#z�AǛM�ǣ�C"o��J������O���EXPTmw*@D�u3h�?P����$)VZ��H�
�FSA�ʅ�Z1�+�\�� �6�W��U=�ЩS����+X�i��oz�[K�'���[n���_���t}�`��Wc�c�R���d!臠�=��ЇhO�:GȈ.H��+_!٠w�{����Xr��{绑'���-�C�yU��E��0���z��+���8�I���Jt�׆[�1h*�*�����mt�P��AH��K�K���Ta�E����Km�es�8��Y���j���By���\������)�2D��LxX����k����<@ԥ�eh�����J�H��n5I�����@_����رc��N�>z�贃q(��8:O@�\��&�Z��ٵE�M$	P/b�c��G�	�
�!λʍ*]���˺��J$�n)����C&�_���c�B�.�M�?����t?��i�\	s��!{�-ɉv�t��<���U%�Wev�Bh�B.�d�B�J�/ Nף��6�t��[���$�
{�d���S��V.C;�Tr���F������"}���8��Y테�.�����~������`���Qr#tW8��m%����/s�Rv`����w=ħ존cH#����oS�!~ڮ]��n�8lFH�7���p<m�~��QR��&_L�FG�@j�(�b~z�J��N$��wgΟ5쬕��؉g�5-�43�ͭ#?����b2u�Ƀy*���v�#뻤�qS68�F��0��A�$��J�fॣ�Q���j��E��RG��Ht�T���9�<�]�k^����2yU�SDx�2��h*�=�� O�eU1�5	ȱ���A63�ynYyuM��|_!k;	8N�X�3��(��O";�qV�.5�/�<6:5�mr���v�l��|�/��#�}�{~���ѱ%��{��n��'?=D½���k�x��~����E�X�M���6"Q�+�q�0������V�{���Gnĉ'���i�����?��?���1Rƻvls��w��Nƒ��Hm�R�:�:q��QǊ�k����I.�zKw�N��/��B�(�K��Be�އ�&M�c>�����I�=A�2����gϟ']J�frr�N��Q�F'蝤Ǘ���+�6n����.�����}�ٸ��,֛/>�♵g��a���g;��b��%��%��X}��kk�@����kpjr^�r�j"H�š�|��d1�jmyY�,s�Z�9{F����g�3f\D?��'�4Umxt���� %�Z͏;�ј�yb|��j�E���Z.+�14<�d�6������E7�tm4�����n���'��6�y@��1	��V�6��?��b�_?����n�R��Z������F�49έC�L������3�B�K�����Kù"��'��q�*C�ȾъWWVhI7V��C	�JJ2l����$ A�=�����Ғ�h�������'[��RF�����;w^�E��ss��-t�S�k��-/`���=XQ	�R��t��k��$P�OW=K�ex�t~j��������������2��<S���Z����oVw~����POU�/5
�z��h���������<��4�- I"]���lZxyi��
tO�@���󪫮�U&<B��O��j�6Q�,*��:[F�V��b��T��a��,s|�*���*�V�z�^��r�y7��2��WWz��J;f�y�M'Vx��I9��nTᗘ���bS�Ӓ��{z_��?�Plv�߉I���逜���@�r��t"�"I1!P��Q�c��������dtgf��^���:�\��'?��?��?�җ�t��AQ���c�]���%E�Ã>(F����45b�E�(i���F`O�D̙։.B�3)Y:NtBX�N����!}:]-��s��O��g:׃6Z�_��_9LG@ϳ��Ç��N���]R��y�ާ��hq�&{O=��!�QL�ѵb�4�65\�K�Uz'���S�o��v�_-�%H2W��S��ߵ|.��Zm�>��&-T�H�@��k���(��Ʌ�+��$�m�}�]XF�HçgO�XP?��d�X��94덍���̮Ծ�o��o1�l��c�`"�0,���W�Y2���ud�9Z�=�	��uh��{iC��/Q����r��J��m�½E�8�h�@j�E��6��C���5b���crH�hyZCݼd ��hˏ��T�˶*h3�n~:ֺ�L�O��-�=����I��IL2�
���1���K�"�?g.p���a�N>�(�rY���𚴶��[���
�w�أvK��2��p2(���9s��w����vZ��f%�u�]7�V�3�ݯ=��G[�/��J����J��駟�[ٷo�5�2�U�v�� ��~�/b cF���i��J�~�X+��n��<�$�tg�0;y����Cm��6⨼�a�Sn�d̝?�K��}�޽;�N�M���Ʃ�c^�j
��r���
�$t�?��O{>�0~�� CO��j��ey��|SQ���U'�]��C��.
J�?��9�n���y!�>bi3�$��J�HS��Ov<�����P�-�J9%G8�	�ҁ��5d���4�4BI]L/J2F"�L�h��������(�\��2	���2Y���ܶ-�I����ܳ���>s�V�U���-����<�أ$F!y��O*bxx���}{`�ODl���/�m���o�v�7�I��P���Âv'~%�2�NM�@��n�>%%�y��x�����0i�������}��YC��E��s��B���1 O
���O�?{�ᝤ�rtZ@�h$��a7Tw#g���!Rd1�mM�f�I��B�p�f�U����Q@�p�D�4��$��3�f���$�ǧM_�ԊoD����Ŕ�����F^�G����n9���6����b(��C�Q����$
&�M�$Ib�,d~�-ϯUH:H��^��Y)?�y.�2z�ja��^�V���U�]����s��8H��Q!#M� �� yԤ�F�l����A������G�_��Fe��D��T�E�][X\,W*���ˠ~q��8��/'�|:6��Y'78<LhW�/BY��t[�E�N�'�8���%�B0~$*Y�����ȟ�Za"6������Ti�:dlK)L��W�J��$PQh��v�p�$��\���w*"�i��S� )�;��V�E%��hf�͖�����i#�_��'�~j�Y&mm�<=0B6�4���\�]�R#��)��SmlNftb�t���\�X���aM�Z�,�a�r�sJ�nY�Ab���2_�0�5Ht���N���$R���?������W��}�~z������s�k�r�Z�g�Z�p��͖k�Y�^#K�	Yv[����C�/L�KDuU��� ���D�E�,B&
Ò���37� �QOz��~�ƃT?i|Q�@jb���m��$��H���&��Ju�����瑵<��a�,�Sm��!�H��*8�J�I��u=��N#�
Ď�$6	�r(�E�=�x+��S����I�v�Jo}Bړ�2�$=���X���ҋ_��@�s�4����R�`�3C+�ʆp&Hec�g>��`��5�yo̿��`���Q���z�7~���I�}�)��?��Gy�k`���G?����7�H���'�$��c�ط��-��'���W����~���}��L����>�/p�S��1z�}��g�!SM���?�+$l����z�ɧH����]��)Л�Y$tRRP�O"w���m��Ӛl��M׹�юw_*��Vض�\�[�C'�}�K�Bb����� �U���T��Τ�hl��W���&'�ku}�L3��B�=�B��U��e������@IĞnʅ:���тgLŊ��3����q�[��}�x���l`@`���3H?)//�ERY���	wHv���T���G����(������֊B��јrWu҉�K�ܹ=���t��wϗ|1��)k�,i�>��V!�@����A��r���m}�H� S�ڕ�Z.�K����:ܷ�ؤ7�nq�Ԧ��Ċ���s?��M}ȩ0xP�-$��{+�Z���AЁ��[�l�H:!fL*���� &)���͗��[�n�7P��?\.�ˌ����Nq�%���VIޜLO�b.[�x�squV����:�$���>��%�����xdη�ǻ�C];&�Y;��_t�.��r����V��ێ���`���E�������_���=5Y��?�ʮߒN��{3���
\��B�uU��׏-�~,�jrݕ��=P�<�Z{�rG��#��G�
���W��p��s����b���l�MR�<I!ljx*8�c�sp&r9�r��N6Ү�.vf{�"m�~�ș�Eݷ/q1��c�:��>�YTĪ1FU2�R����>&ex>OH�ɡh�Z�%2�����u�J*��1̠�AW]��A�_��iTTs����Au9�����{ma����^�!��3���޻��Nb}����暷�گ�x���� K�FJ!���|���[[͖�����E��yi�j۪Ҟv{R+d�H�nl�=�����r��)��������a|��<yrm�|�����G��H��ۨT1_lm��	yn���v���x���C0bۀ=�\u=@�H�7�e����Wؓ�I:�J�˲
ج�ňHJ��`mC�6�%y�D��Sx��Q3 ��	��)�_���"��3B�N"����Ô�˴�f� wx�Vc�*g��P"Q���,���z3�=��i�-�9��A-��9���m۶)��2��V�,�͐A)�1��@�P�Xz��C��FU�{�k�+k+q������r����H~��N������Sd��}e�ò2�##���KJ���
��Yz��1	7p���M��� �M8��3�����(�WS�4�J�I:Й�֐Qhp��
�&��*W�jЉeQ�%'wv�sDY�"��������e��/�V��]"�*�˕2x�I�]!����Q)J��`iy}cv~�� ��ϣc~Qk5�M�%��Z���~+��H �Fr�ի@%1�����d�ePmF*���4['L�XN�c0-y����HYYo��yQ���4Q;��F��iG	[��t���~��'''E��S!��I"k�.+2C���9�A`NQ�ۉl�mo�*Ο+I�6qQ���O�-.�~2�\�du�+j�aA��B`B|��^�Kѝc�M�}�m��G�-|�s}�;RD�s�q����^���go����N����7c�m�Ni��C��w�)�\�c`kUѵ����g:,��QW�mE�x�p�T��j�s
P�C�^T#p�qL(ޫ�Ny��,�I��N�$���G�NrTW�tS��?��ny�-�`����ZB w�yg��G��sy4c{����%w.��vĤӰ�S�["�C?$���%���/��1M�E?$ u��7�]>|����o�Dt�k��':><LǦ�A�j�w�񇟿��b�����=qɦs��	��R�w�~���S��vRĪ���$���cAV�1�s��<�3@�˜ 2�y�ې�v��@p@�h��˅ȵ'h
QJOX �+xDL%��^ܝy 8��+)t� ��z��Y�PltS�M>�d59i��N`��b� VQ�Q�e��F7R^E�M�k�EިYG9͹ ���'�j��i������+��M���������K��'\�)x~��<0�'�*"�&�YWt���ȍ����B�>�pAK�sy�î|��w��t)�[��KB�Na�q�Ų�y�O����h�����p���j��0TT� H�o�'�F��z��E�-����'��
����v�z�_�g���	�~��%:J~y�{�'���$Y��� ��iϚ�����D8�B��B��?�0}#Ɖ��6��(��y�}vN=�c�EW��~�\#,��挑^u����9�L�9?�9v��:�@��5f����H!��S�����ݲl$��έ\�F�b�T[nݰF�d��t���r��b6]_S{h�8ǔ�1	K��=��-��vUy7�}�Ƥ����Dr����n��؈-�(�NDo��b&0ҟw�4�"��E�s����k5V�	Ƒ:(:�q�zF�[Y5�-C)�Xa+��N;�H�jkk��oz����g~�Go��&#�Im`h���o���Ȳ/��ɱ��;������ϒwO�4�,�͋�Ǵ'��2O��
t1�59�t��t+�ڬ���?��?&����!Q�z��N������69��Q�l�h3!������ι��(��\�\ͥ��©(�N��QWÖ�+-N���|4pC}�~�Pݯ2�^-2��L��L�Oe��k�bNw��hT�ldr$��HT%��T	��ǆ�R��.�Rr�U�X�uE!
**)�$.X�d�j��Z�|?q]�⠑���FG´lB��/���6ÍJ���-/pk0 ��2yFU���b�Y[OcMJ��9�jֱ�8��00�&,WV�
��n��I:���K����S���4��Chs#�G��	����3g�����Լn0�-�� (�vT�$��p�t�O�i�	������bҒ��がF�nJ͠�ϱ��֜b.hz\D�I�޼��H�AZ_ѥ���v�'%��c�!�ܧ����o�s+`',���Az���3d�#�^4\Pv�����R�NM������M�(�t6m�'e�K�Z�.-{cc�c��01z�br�5C7|9&�	�F�6rs	!'9U���{����c)I��S�>�9�iOiךV���;Df�ÈsΫH���n�^��e�]�{�nz7B+\�G7���RZʜ91�9��~��� A�� R�����z����i�O9�7�G[J��E���}9(;9J���)��m�����s�С�n��>�Tp�W��p�P�8�4ٔ�Tꂔ��.b.�&k��/!*�z�K�y��^�ߣ��C�Ez���&澻.k#!߾1�~"g��ID�!a�/��x���(*mL@��z��	��
��[��57�ʓ��������v���1m���*y�+���.�eNS���zԐQ_߀�������^tG,pG��"��"���'0I������u�J�Bx֙k3���^��+���7	�@W��Ojel�}'8F�t
���b|�'��1;Ί�7b�%� �QC����~���}B�$Kz�d�͘$�VCH1��]��
8DA�Ve��9y�ȇhL
�k51�Xv��������	�]�c#��~�i�R+��_N���(��! [K��}���S��CGF
 �6|w�� c@��TJ d5�f��,�����S��+<��K�tZF5��Ȉ��$9a�K;�~��qt��K�8s&N#�.3�f���C�˛l���x ����c�L�ݤ;/���&	�u��*	zC�D�ad�n&���	�������l�5EE+X�Sv���s��UZ�E2YT�\��s/*�t��ER�NC��� �6���p� e����g�%�cٺ�]n�U��s�B�s�3 �씘g�����ER]ܷ�0 �r�Ɠ�'�E2����X(�{�w�G덓sH��pf��RK\_�u���#�U�:���Nb_����
���}���T?6��Uą�n���^a���ϯ�6�f�OM��ܹ�Ϟ\[^2P�P�[I ��L!�uuv�T���Z�~��WY��.
Y\��{�>i'u����7�]��jV7���)�D��8Rx5��z&�R?�ch�A j(j��r%��А����]v��	��h}E���j�"++g_������V^�ŕ�L!��Qmq5���~�؉O����?�q]3�0��/|�_���&&i�
94|�\�T	
�/���y/ qfR��$w���$�+�;z��>��?��?'�Du���(_�� ��R��U�B���7�084t�����o-8���w�9BO=��M)В]���z�������l$t�D .Ry�D���hڞ�&����ܠ� S$�D�'s㒬s�����ޢ�~�-Q�r\n�a�2,%FU��LƱ�	<Gҏ�(�
S��erY�U��=_��5����o�z�'
g3I�=����rMLp�����e<E�x���w�/ȍ��@�e��f=�ܙ���*I�Z"6��|���������d*�`"�Z�y��뀴y]��"��K4�3������v�=ԅ:rO�˕"P���%��%��.� �,&�IN�����/%�|VU��4ȦN =�t���IV���/|h�E�?QD��M0'w�݆%#�s%�nC�:N���C�nef����3u���(�.�(kyhY��0gg�JR��.���У�]�7@�/�ܿ���W��:wrFZ^>qf���*���j���#�;��%��7�88�4j�;��b[Y^�SIZ�����F��g�,�x6���e���k�e*&�y�w��E`Gh%)�Ph_�n��Dss㇔���t���K�ĘS�+O��̠#,��Q/�U��l:�Idi�o�Olr&:]�*^�m ��
zj�M�r$��z�N��Ʊ����E�fd��jHM15	��TĔ�C�1u���O;I�v������^bz����m��Q���{�K{/�EP,��EH��-�Ź#4t��(�,.$��b� �ΛR����_}+�����"?���xX�(m����-���;55����ͣJ�G?��3�<�;�M�����{Ag����wd
��T~y����e-q(�2 &Hא�X\�'�OJ������>�����_%�}�vR1�;p��W�;{���|z��n���^<��SO	�|����o���d~���Ѓ�"�L���x���n �A�MT�h�յ�b&��;�-����[�����G�8�+<���i �Yl�����w�r��}p�/`qT����Cw�@�M��]!ole����I;��!�a.��u�]��g�-3���tA��`�$��Ag����X>1qx]BUt��o$�-��ق܏��EU�ԉs*|tBz}f��}9CfA���$�}��k{����3�uK!sI�p��H���O�h/P#��� \���FJ���n[\3fPLG�6�L�9q"��$���6f�7LjL� LT��@��I2�R�.��{ͼ�LuĦ0NUM��װ2�?�<	3�U����]���.=u�$���4��]S�t6��A����m��vaq��}?{���[Q���lt	ާ�I���<���m�ܹ��kҹ0l��g�>wna����S�����j(�r�0���y*�1lZ7�J��J�5�f�Q����屝(s�7Ch�Q2��$�'��+�^(劄M�,��_4�|GeJ�I��(`��|�y��E!�;�m�&�/�})e�J�wF�q-�&��� �hXz����+�j�[�<��7+�NNR�-���e�I�]���b-���M��Lvlx8��ӧO�y��:�j�Irl�����Xo��.b��r�]u�)��5�'I�6CH*����fY6��6*���a�5۴��7}�q���ىL���5I�i�[*f�(��a-�j#������l4Җ��s`���GԤ�w=u���_�5����6cǓv~T�$y�ջ�$��7%x���z��k�;|�p&6����7�t3!hR�	��$)岟���	"0^��J��pp����4
�P�^��C����cD�M�0�Q��)&�#�NZQ�@	e��Gra֡Cϼ�7~1�Qx�+F������w���O=�e����d����^8��~�N�!��Ҋϟ_�0�w��yǯܸg�?����o�;??+�̵&�M5��Vp���t��ê$��D���\��䗒�L�e5�����ź���M7k�=-U���YI����!���جȏ2�M2���&O:��Z�4��۶]�gdϞ=�L����3t�3�^$����>'�>?7O�Q�����=s2;X��9?666�̉cuя���\��̬���u�}�v�w�dv4<��]~����KKǎs���>���������2>TS�Q�{eyUo"����B��nH�C{��u�P.��fщMrKc�o����x�¹b����Mw�E�����ðY`��U����T�Ok幘ak�f�o
���G	� uwJYI�ZYU�J�VTQ�*dk5uP��JK�%=R����R���3���
�|)��b�p�Z�\L�M-�����*��}��U�Z��j�FS���{��T&{`�/�bZ�##k��>S;Q�~|�Lf�o��5���ןV�#�oY~�l�9@��)�vz���u�$�Z�ջGL�v�� O���i{`����J�L���{����=[l��Å������w�J�?=9E�37�B1�K��[���k���GydƏ�k��y��o� @㹮�a��ǎ����N��cK7邻�@�3
�Ez3����/�JO��y�������<�K��f}};���J�Y&�JEe��Ɋ	0t�[C��'�=�庫;���N�y���Y�%[���-�En�@�!���@�]�6ɇe��?�,	�!���!�1ƀ.�WIV�U������M/wn�������l��1��yw��_;�{��P&�!�&&'���J*�)*�E�@T�ڤ��,>5��ҕ@p��=�/�E���u�>�Մ�"[�!��ovw�*�=8�I���2�[49b8�0TR����1�����:Ǻ*Q�pևӨ�ӟ��x礔#���y����	 ���|�q��ؾ}���k3Q���]q�m�}��_=v�`���(&��r}�i¯�ݦo7`�
%x��s��gM#C0^ev���,F��Ї>�ߟ�*\|�Ř�S�������0L���
)ߟ����������첋 ��ځs��K~G��2�N�h;��\r�-�Bn������[�'������0�#�^�ϓ��0��Tɑ�R���T ���)A�ɾ�/gD�='�Eu�*E� 6 �1j :�����u�b���Q��<���a���*Hl�f����$.Q�xag������N�<	+*3H\����J]Ո {�t��a'J�����{Û?Iǜ���C#K�Ή�jˏ����t�"6�GX�X\ u�F�ܲ���ɀSn����9�R�qhDAO�۪�ed�B���+K�����d�9y��m)g��NM��^�y/�61VՅ��Z�^z饷}�S4�
!�S���9��n:��s���/���k���m���'s�x�������J�0*JOD�-�׎,e$jp�:~����U3�v�����N�_�j��͛�-�&� ���.��C���3lٲ�x~/Q�u���+�����������G>r�Wbn�T�q�E�mb̜\����x㍏�<�Y�	ss���Z��?�S?g��Mfg���ʔI����8��,�r�(GB��m=���.~���z5i,�fڵ��~�� ��D9m �uHd��P�V��I�D��1E�Y��07wlt�����]�cQ�,�/ t� Z,:<<\�9�Z�fO�68����ZyO�J
��~��$E��c��9���Qْ�+B�� եR���H�^|�P�ur]�5����B����׺nju7�e�n�<b7�4�Z-ݶm)�+�ʵ��w��+W��?��LWDWn����a���7�*�����ك��gf�0�]��~b��᷹��
x����)���.No���%�\sM�H�O|��7���_������0ֱ��������]u�U�sy�.��S�e�n{��.��U��5-�LT*�R� �'7���p��y �ȍŎ���"�L8(4�OR"��r�<��$nD1 uMŀ�Vɕ\�x(��dE�v�Z�r[�>�Ti�����
����{߽��ǣ]]ӓ�!V�:�K@p��V���x�پ����g�g�)q%�� Y�f?!Ѡ���f:����j�5FI;j�J<<���ʕ���L*�Pכ�CUx �X��u�7��ʓ�v�R�*��`W:�깙;v,^6rt���K�hD�ӕ�]v��sɅ�֟��sP����Y9|�#O��Z��g��[�f���W\vdt����r�wdxvi�<�R@�U�a#+!�X�8sE@5�&oL�X�����}���{I��;Ԩ��N�\b�1  ��IDATL&ׯ_�uWa0�-a��)������������������=o���>��>�߯�}�o*���������1*t�vECr���ģ���㙉$V�fٳ�9I�R�$d�iX+�-��}�gq��/�p�y��Ek�Q�FFÙ$U�B�OOO����o�ihO>�d]61�3��l�o�cۙ��tx��@�����|ц�׬J�̈!��wd;���� G@��s�Qa5v�������~�_�+ە�y��("��<<��s>��y��e��0��)����a��#��υs�б淰Lo��j�'-�?���,̊�;;W��
5<.&�Q̳�����I*
�����:�Qp�X"�{:�"Ј!�/Ҋզ�{O��Y��Ak;2n��!���Ŕ5!��1�)�S"�AC�Q�e�!�.�V�VL��Maj2�-�}C�F>��B��Y�eX������:~Q���E���_���ݍ��V��k�;��U�������SO���� қwc8�v�����eV���n@iq����_9���׾q3�#c�c��֭ÕD��y�kP� �+V���[0�J�k�����K/a� G &�m�ELg���'$�޻w�g���$�o�o.�;x���͘™��O�����y<?�6-t��nD�;JB��0U'>	�o��(ƀq?�S�/!�k6	��Z�8����.���7n|��WcA�� �1�(�!�V�H1!M"����������i&�,IR�r�.2����+������C����o�,{͚5�j	\<� tQ?���1��������261��r�AJ�
u�I<�[�n��b[�B��a 	�<��sd�htR�KӸG����%樅i�[���f��!���NSG����p� Syv�Щ};�a��6mڄ]��W�W0/����ο|��_ dd�ʣ����o~�'�]�뜸��(��2��&,�T���!�hz�ݏS�i9p� ��믇����@.7P��}qxV�Ir֦��	�{Vd�����;�v#�]��aV�}	+r�_~�Ů�T*	S�:��@��d'e`�S03^t1~y��@�.��ϝ�1s��kIxQ�''Eс1�t�W�^�q��`�p�-�x���Se�(I���l-|�6k�R��U��aU�gyT%��S��,��<g�`��:6Y�X��D:M�E��Y7�(�2N%��U�V�?�P5ig�NEO.��1$:����,��3������͒Y�h6����=�=���!&\�;�+���?���#z2�D�a�s}]�b	�l#��!wtI~&�ߕ��m~`��tL�O�ؾ��V�x�mU �q����Y�}�Q>T'��>��#W\vqowfj���}�݇-˵���3�J�;���/���f�r]n�㴹J����k�\�ìە�_Q$�����,��}Yz��m��S�}Hj�������M����SV��Y���C�N$�zd 9v䍅�hQ��pj�CYCr�n�TR�r�\/��%����H|%5,͓䘧X��A`j���rͳ��G����)R*�-�ض�l$!����"�\Q���p�)'뢸9B�Yɔ��;�e#�p�����,�����æ���<r%U�������[�����gK�
��ԩ8�o��&DN���)������@Tt]�`3#�)0uWo��?��G����잟������#�����x�)�����H�S`g�/_���ɩV�����/��|�r׮�_:01���)�7|�ߔ��yk�$Y��5b�H��jQ��\�_�Jz"�s�|~��Uz�R�)N���-k�� �ɪ]�љ��R��_����IdcrY�}���U箾��t&��ˎ�T'&���8EejE��XR:<z�;�#�J6��|�;#����n˿��O�Ń�����7������C������y�Lj/�0�I,�:1"��Ty��%��s9���(�fL2p�k�T���>�b�������ʦ�1_�]�<A"K�ME�J�r��\�611�Mh��2'�n�����P3�:��)Y���ݯ�z˵�x�r6>�LQgPˮ� �J$�A�e2�L���~g~�x~|t�H���T��:�5g�2�"{'Eg�\��1�*ɂ1�/�:u
jB�ۮR)`>t�H�cӸ��ѣd�%\�=�:�z�P�׶W(SBM�.e�O�ıȉV�w�s�ps����,qv?=?�#����G�;*��.�l��	hQ�jC�҉|m&�Ȉ��@@d�s��wv�V��n�nh�A&��R�>�W���n�(d�\���E��$�L�-pɷ�z	,A�+ e|�n�=$�(�,_L,�C��\+T)� ��;�\`�����@[�}�]�G`���_޹��_x�{�W�<�xPX_����@S��b6r[B�Y�����[|^��.oxUJ�(y�=�`t��c���?�����N=v����.T��
PO���ۻw/K%��ˮ��92S�X槧qg+E;��m��K͇fB���^�Y(�5���4ʘ�9��g�Q��OhQ2A��d��� �Y��,z ����(X/���`W�~�V�Mr,\g�B��Q�xd��5jc)� ��(��,Y��ee�����>�[��t�B�*|�!�q*ǝOB�X��#�`�����IK�g;��*�2L@uE?!G���ȯ?	��-Jd�v;��g?�B�z��.L>�\,�W�^}ᅧ�"��į�wP���B#v��b7b��{7�?H(��$�kȢy�d�t��ۧ0�T6�����h_�����(w��x�|�$��
Z0��`I������$X]z��'���*=�е�^ە"3��?�)1�Œ��<�Ji*U�@iS�Pْ�$Q��q!�q�7�8�dʔ��0���}W�P�G\�O>��Z��O�ì�]�X��I@�Ԇ�c`1�x���
8 i�x-,�/�������*$��I�vq���=��g<^%�"�n��W�\�Y,���ۋ�/Xc�K�t�}�
�&,0Er�#`��Yr��������g\l[��CSY�z;'�`���:>1sj|j�t�X���=w�B�'�n
��N��Bm��x�*K(�nrI�\5��d�\����j���;ř��}�Rdf�&E\Jgb����%��Ĥ��Z�� p�q��TJ�B
6VD�j�bF����MI���ڎN05pj��F9m42��PWϝw~p�L��'ƎC(�������������G���Ύ��~zvv��o<|���/�ȴ�;w�8r��<p��!�
�."��t�ep��LK%��VG��,k�����^��ޑ�x2x&q����������.�c�N��!����I��~����,�����-7_q�?�ɽ���:�Z)F|���.<g��>��s�O<q��?wӽ���zŷĸ�M�i��{Vf��d�MI�G$�0(��Z.9+fF�1S�	By���t��m��s\�as��@�t6��K�P?)��<ei����<�WW&���㬕��D�_X*�q��ȌQ�R��\/��C�a�lQOsI�.�)��v�<�[A ��T���NG:.�t�f;�-[ֿ���Sc^= +��ɤ;��x�0?4�q�zNݵk���o׳�Hya&�xV��Z�З1#A=�׮�b�`w2�:3��9�<���l��G>�;�U��ѽx�}�N�>E�y��=80�Z��d�t_FI)zV/Z����[�� ���{i�KX�[�nq����=˅ ��T��34���~nfnj�
�aW)J�?85?��Qt�#�*ݽݿ{�	��x������ܻ�R�`�v��v��s�������I���r@Uoe_[�5���Zܬ�}�x��g"Ɍ��6�:,I p�K"��^CY�zզ�6`���N	yx�jb���C(��kH�������xZY�;V��Jy)�p�([ Bl���zǏ�FT���Cmwv�%�Gqݯ۰�)m�Ti7SX�n���SY���PwǢ~���V�V�E����jr�Z��l�ن�)B�V��0 `R���R�|��/�J�Da�<ׂ�?1���6�<�K�����gD-.��}"���cEbC��X�2ӌ���\j�To�Џg�E9io_!5k�����R�*w�mq�g�%g��ϒe����Z��a���W��5Jb�����К@#j�<�m%SqgTʣO��ok�}eB�DA䢫a� ��~����,�"���'�,���Gk׬�w����p����߇���~����P(1a.fQ��_���r�rp�;&�=Q���%���3�6�d�����ǳ�0>�ar��o������ql�#oS��[o��'�Տ+K�S�͆�)+.��-���G>rӔ-����藽yzN`4M@+��4f��S��P�s�5����\Etr�����TZE��`5G;�;[ uSn��"�=��}���5�i*����?kQȪJL;8eرl�@���2B���/ ]�B�z&��n���Gf�Ⱦ#a���{L3�uvnF��$���&��J��}�p��ujv�[&��0� ק���x���|�3��/|�x�끘fS���%)��cMq�(R�Q�yڤr�k�r�=s�*�k�x��X+V��Ws�&}" wtݺu�)<ix���E��+�J+58�x�]�vmߴiӒUK0�}|
��k��?g���>��O�}��8&x�E"H�P�#	P�;��Ç%#5�re�BY:���yx��W�9gD����R ��7CIlq(ϱUQ3���E�"����B�^g(Fƺib�pƱ���r��H�m�V��[�����x����(yqp� ̮^����]��~�}���b�g�JQp�s72~�[Es-�R$�ڴX |���G�`������M��K��Q�7I{�$H&�z �pCạ�����8ڽk_gGO,N�葘A<�[�Z���-�M,�lwGM#+:T4��Q���nr7��c�S����oզ�ǩ�tU��#��a.wE$���R{b!�>y����U�2]]�rJU���R&�kd��f�A�{'g�����B�T����ް+99��_�k�W/ώ��c�����a�x��#�x��犥�0i�X�;
��-[�\v�EK/�`���?�������De��d:xyAC�̂�����T��y8���ˑ0�=8{�uY,=��X/���;B8\y�s�mF�`��#
_�
�vۭ7<p�[oݶm�#�<���q�۲�~��j�8��n���o �q���ښE�]|�C?"NYo�Z(�kj1N��z���LgO�>ח���=A� f�r�,�ac���\!W�U�z��15խz5�&$[�\���z��}dI�DQGǑ<Jp�ԃ%	}[����H�f���Ӆ�U�t��R1��1Y0.�s���@	����d*����� ��vd8 ���AE�J*Mez��{ ��-�o?❷f������l��OU�z���/d�D�ި7R����cٮ�x:q|l|��PE�f���t�49_T����쉛�{ V�;��ԭ[�b9܆[��������n;�ﭱ�r`��ټU�f�(RMGG��� �q��]�#���W�f�X/�R�Z%�;�}�ʥ�l�2�����_>_��\�裏.9����/���v̰U������'��3��:�m�^y�_����r�_��W!�8��믻�ر�k�=�я��1<xՕ[~���D��,"IQ�[�\.]� >5vJ�d;:s��|,�)���y<��|�a��=��Y�7l:��z����!����U�:gO�T�@��6F�艓��U�m��pN�ɊJ����A�Z�$p��|>��(�<569�z�s��#W_��.B�٬�E��)��.�Ձneyv�O�d�,�oE�9�@�ZNv���?����qX��&���A
@C�,��D&����[��&�V� ��Lf[!D��g���T�{�B��s�=��0L|i����
��p�U�g�y�������|�J�\��������4X��Ud�������M�e�CC��sud����kC��i<	��������agc���S�G1F&� ���E�J{��<�7�{����W�u�]Ў6l=z �1�;�3�J�]���c�lp'��]�Ps�
�>�~��4��h4(����T��V�ck���6# |1�S�Y-� ���/��Mr��W\��SO�O���]���[�q]s���ׯo�M|*����[�Z�g��O�$|����8.M�n�?�gI�i��Zi�g-�%?OGg��G[d�d�9.ǥȄҢLC"�΋���Z�&kC.�r�kb��1�/<�,���%��"II0��IgJgqX���]�l:���9఩�9a�Sk���ȇ�{��˨���&�
$��͆[�JU\�j�"�
T��X���o�)�?�0��N�<��Q-�@����r8�HQ��#`4�9Y!#)]F�H��L<�AjB��s�K8:N&Ĝc1'�Bp�H5��}�6�bf~�2h�o�������!�_���S��KVS��e���~�����a�力�oݺ��m�)��'B���B4�������n����3G^n��$T�X�-��%���/_�W)�%k�ѐUe.��9u
�o�����da��m��?_�r��Ȁ��#σ_1̉����`;��Y-UJ��c�Ϝ��@è�Jc��j�^���1jvF�SD�	����MO������j>f�p|/�P��T
3���X��7�k	�n�|����K�!��������f���F�yYA][u�>26m�q=�bE�U�N�(�]W/�j��"l_"�Yé�%|���˾�P1��^�kX��K�����88�VVR��:Kf5�ƭzL�D�1�r�ֈ������W7��y9������nT��VV})�Wg�P76�p��v��j�P����؎�^�zC���:2����?��g����;���X�<x譁���c'/��mqm7�HaJE?B
���-�*���MZZ)
\���X�K�Ё�&�n�ٹ��ס��m���}y
P�X<p��N�Ί�׭]~�]?|��W����D+j�޻�k������!�zwn�vߏ�)Z�@6Q9}<�����`�s e�k^<���J�8�$K�AU#�Lߥ�S����:��P%QhS�(��V��r��X��&�^����4!@=3)hKdٶ*�HT<��aU	����'��2��H�*�z�X���ڹgo�F����xRV
i ��+6�C��!D��Ģ�j&)����fP<&�Ǧ��<����s���V�N=��7K%�WO���H�ſ���}��_���zv���l�3��E;�N����I�T�zh6;,�^4�Y���e"y�2E
�_t�֣'���T��S�569������4pb������-]���)�AՐ|*m��6;�a�5=�T�\C�����r�����C7a�S��g�<�/~�v����j���O=��9��o���6QG��O_}��_9u��ݿ^��+;����g?�Y%����R�!�O�-{f!�)M$)
�M49���NJ/˪g���k�ҝ���I��9��>�l�ߗ�D��&J�,1u�1v��^��T�������=Ԁ�w}�6���Re���)�T��8=Iv��� 1���ҷ�j��R:��H��J�#q`��k.��i����c�gsL�K���"Sh�-�v-q�	_���X���<��$��?�8>��iTl-:�>|

�WB�s4>֎�4Lnqh�g[|/g�aA�ug�X�<Bb.��Ū��&?�xB2/�6*>E����p6<J!�e�3R�"3�y����;�Ë���dA�:Tne�H�Lb\��ӓ���X^�d)�J���9N^T�x�|�U,��Q�$G�Q`��#oAX�$�ݻws�Uog`

w�`�z����>������f-�qM�����G, p:�����O�D,���.l�p��g�\��g��p_�M٘��ˌ5�9:m�.�������M��V{p:)v�7���/��\c������#�j@��o�R��s�c�Xzѧ,���(.���D��zT%�ą�RiK���{zzZ$J7�e����/<�J<ֻ0Uz�h�_)*��tѧ>�9�մ�TruFE	O�A��.8�)����q<�|$�V&	4�ё�J	:�x�6U�;��	'�?��1ܺ�$�S/S���u�0W�Y��z�adV]����|��f��/v�'03�$�;w�Kg;��Յ��G�իW���E�,L��C���N�����/�SON�DW���jˇ�FFF������G�5h5��*Q>_O%�%�� /�zD�j�x�2�"��hVPe/ɱ�C�]�S}��
u��@�B� kxfn�:+����o���,�n~�[�Z�fMIR����6��H���(�AD1���	��f��67 �:G��	a���	����CcO��#�����N�F�+�`-���޷o_��u�Qs��*�N���>�9��$�����|��'q�{�*�-N|���~������ڵ����];�ȵ�Єdb n0V���&e�4LA ʋ$��UE �?��r�_��s{�q܇��i�-�핉�E
��
?�Dv*����}��SH[inn���b�T�⳱8���I8x�b�Б[�1�=Kt��U��KM�I��ԭ�se莸$TJ��;%5D�g� �K��ծ*Zl0���d�p�^6���|I�#F\959d�7�X���+eW��_@r2�l�Vǹ-���/u�Xs�e���{;�o��T�?�p	@²
�ʳ/��x�JH|Yn��g�+�����}�)��;�?���lق}v��vd{�_*�����v5��/�lb�xhE�
��v����ʼ7ђ�k��`F�����|�%ڞ��Ý��������_���������Ԙjw~�C$"����c��������=����|��z��ڵk7m��f(���|w���Zi��eبF�b��L,�B���Wgωl�j�.V��%dM~tM��e��U���x�6�D�\�e��e�(p��z��\@���$M"��m؍jmnN�+�\ �[��?p�s�Q�����%��E�?3{�3�=%��l>�la���7�/�K��g��O����>�c�ɀ�ْ0�@q�$tŋ;���\����,���cR�33�6���E���	#a-%�i ������w$��H�Dϼ��0DR�Ql�� s�Z���k�J���>#W��!� J������39&F�2gl����R��B�hQtz����j"g?Q	�j`F�H�%�q52:zb�����dlE;��w�KQ\_�*:gd)��`Yf�o��ï�|+"BٺF{��oxrrrf�r��X�a9P��Lw�V�_"I.OBLa������rPyk���Ͻ|�7��k�bV���4Eq�rRY�M��p5�<����>"�{�=��F<��q��ŷTe[�Vs���g��亩����W/ߴ�ܑ83ID֑t�����ˮ7�"�|�_�L�dG�qb���h�T��i�*-�����2���T�Q��Q�{5f_��b2qYs2!>�a@\y��O1�
���C_
��VIjZ���l_ҡ�"�u-r�z�Mb�צ#�0s��q�-B�DE��� �Dk4_�؆ ?f�eM��	��W��?��������Y��&�ӉeӪT��슅0Y���>7G���lP`P�l������ݍ:5Mܶ�W\�k��0��?��?�~��Y�u�����G?�f��{V���X�VP"��Ɖ	B����u�!��y&Gn(i
([t�0��3�@�ٜP˝��V}rx��X��m�f���m�51�O��sƝ���o��/��/��|�/���#G�`��ر
g���$Fq�'?�ve�֭[��Q����Q�Qꔱ�^TY��M�ǣM7��E�!Ed�D^�h9,#5��ļ���nw�De�����3�bJ�̊#D�s�J��?9)��$v�U$J���M�(W)߿�x�e.�)���K-Vђxi�irll���������e�����\��EC�J+�w�ޥ]��b&��h�B��"	hH[t�Cma=�,hB�L�ZW�D/�.2�Ƞ�������-rɈ���41�e۶m4
����g�1:�J�D��H������#
U���1�-�C�����`�0WI�$n�����	���A�3���/��GF��F-�)G�$$�r�:�ȼP�����j�� ��D�ge�v��������*�72���v\p����_<q�}��ҪU�F�
酣Un���Z92���<���7��o���_>��(�=�,'|5v{$�;l֓���o�q�4�O�&�� *"��{"���c�0`F)������-�M;�!�$�cJu���E'�p��>�Z�%�jS㱱�:k .���k�,i���	�Y�U�@�Yc8�w�sA�3��@��B�Q�9�E��&�@��4)��_iQJ�X�]�+-j��ro�wK�@������u��Y�N��ٮKe�����D&kF�j�ԑ��
b��in`�M���38�3��~��I:�Gy�Rm�0?6>1<��\k|���p�2�W^y9����?Z4����˵]A���>�OOB&j��M髾��f	�o�aG'/�vg�},�:wDa�~�r�X��*�fW��^�ߦ ���Y3_)���,9v��y�&&p81������������r�|�<95Mu��/~���(ףּ�];u�C��lcթ�+ҝ�mz�??}���#�;�Xߐ S��@�8�J�u졸��z<b���J�[�^z�j	"��R����<d�!����S`�]�A@���3��r�͘��퇈�ͨ/+� ������[��GRC##�]KHK7�("Ҥ�Z�^�pv�rX�=�T&R*�D�X�`����g��:����ł'���S��~s<-�¢-[M�X�|ir!�QLU59�uɦ�:�t�˦"�BŒ�t�p�V���T$7�9���\.nF\Ywe;]W4[�L5���<9���Mq�x{FΤ���2<Br��%̨S*�qŲ�
�9�"��K�*Q�W	|���R���9�1ų��<P����I��e?M�z,��c%�L��mձ��R�QW5쓜U�����ҝ/q*'ƨ-�`����]4�J2�-�$)!q���N��:�E�Be�P�ec%�����{�,��@L�,]�����|�2��_?��>��m���e+W��a �Lķ!R��Om*� �	��cs�s�mh�Z����n�������%�bjj��0��s*W{c���8p��a�{���@_&]n���R˗*�8m�Z�ls�-������@Ir�?�������;LEg觵
٤���th�s�R�:�m
��L_���#|�>9��y��f'�����~ۦ�X"Ϡ/�Da��f <W��l�;C�Ϻ0,2�[e<�P8����|���S��g"�(#Re���e*jnE��8p��u�XAe!��=A�ƴ\K�
����xr�z��[�~������#�\��Z���4� ��;�3� k���/��ˀ���1���	P:I=}��>���;�b8�q%����z�8���@�x�t�[P+�63�����y�xo4}��5r	��������)r�$ ����z������?����?A�����M&��#2��`l�vw�`���Ox�k���&��i����OO��#'_)7]�Κ�P�Mt�2��1sI��SlR�s��k�e�rM�O�[a�8�s��%><2��Ll�[@��,��:M�A�e���'�^q�p�)}�@3n2�-e�E��x�N�xC"YR��E��(��33H��gx��=�\�+��F��I�dA�_�I"�A����-��Dl\9�@�*U��O��`:N�	�e�El��t�MCd�bY�<l��i|�9jDe�;+��^ˢ�5���,�J�]K�����T�߻x�ۆh�M��ѣ�dG�R�b�Tw/�$_*��WKһ�u@~F(9%:SecY|
C��1�?�p$��^�zv,��ԙ�Y���k��_#+G��46�[�v�,�͘e6�@C�^�Űs��ݯ��aÆ��L���혟W���>�PO��W����<�
oEU��r�>�p����ȭ�A[�X(��On�W��av�*�U�`f@86+�Jf�Ƞ�*�%}�+���~w,��F���^*�;o͗���/��R�N��Z<�>6u"�bT#�P��T;��z$�5�ȥ���X�j��$�9��J>�}��-�*�Z��G�h*;�+�{��8�`J�����R��В�2 ���R1� ����JW�E���:�Fš���R#؁�4�<���٥Fc�S'q�q3���:]�*1Ř��ܾ�Uϥ�,3#�KSw~�&/(L?M�(�:uꔩ��|�ų���B�Z��ܰ���f5B��Z�ʉT��-�u 嘱�9�z"����Z/l �赺-���04.������'�C>t!�9���3�����r3/�K�$Y>C���ް��N<���|��~���g�*�k�%C�3s�����l�^�����Wnߺ���k������S����/����Vf���Ԑ���D�|��JB4vo���ȵ�E�Rw�@eP�z4�q%�������:"^��?�Q�g��K����7��ӛJ���XR�u�y"�NL�d�P+D21M�R�HB� ��B
ĩ�q<��\:"7���Kq�*�'�|��������)j!��f�f��ѕ����Q�X�Owu�ҥ����b�+���F�dùJ�3���ے�󵄑�;~���m[W��h���dOg*1�]�j��m2��s���f�̈́K6u�kW��$w��1<Uŗ��HD(>�������x�+ȴ���0fzc�iϗu#a�,�nLU����wj�\�Q+�Q�2_�'��&���$j����l&�Z ��F�F�cu �z2��l�����tQ�$�`DZ�[=���Iݽ�khH��)�4�����&��Ι�o��oR��Z |�$�JBaƊ�z���)q%���j��Ǟޕyc��ϕ`�e�.J.���X��K�j2���E4�%>�ւqJ	v��lb��ps��(�g�[����9��}�ٱ�{I�c�e˚�T`?�<�}SR�3��3.�34
��W�X!����0~�WXo�·����YL/�Ō�۽+�kC��H�+��袋 z�����p�Ebߞ_(G:��'O
G��V��f��ϚU��HS��0�+!>"D�ފ��)v�O�/(�L,�����ʩQ�({�78���K�f4��B]�H���\�h�I�*�'�<��L�b�'��OǢf2�~��7�C���T}���ė��B�#@�=��=��w�-��xC���'?���{9S��#��7˧���#+�袅'g��+����	��"T �,�S���)��%�9e���F�t��b��V:<��^���_u��{	�400�!��Y�v�@��/���������+E� %����`n_w�u�v�J���K���F����e��n�b��)2�E��U���H�"E�;(�%jP|K�:�@؁�x�'F�J�o�g�-&
���p�j�[r��RPU1��.�ЪM�(�kF`���x"~'ץ<��,�1ѳ�	}�����I��[��&�O�����[���>�i{bϋ�y��N ���h>۞����B��w�Zp߮��a-���ZJV���
ݝ�ĚU'K�x �&�R�oi2��`�q��CV��H����T�{��R�'&0��"M+Y%���9q��Z���]��ϾJJ�� ;mb�ڦ�����}���ޝ;�.%�Z�I�Q����={c���0a�!�L���=\}�Y��N�x�/������ !{�9�B`Z��"vd��<e6<
�ψ��Z&���CjR������=K|�2�3z��K(G�*��\m�P�˲��z-��/�`�c{�T,b(X!�Q��J�V745�M,
����02�aU|��-��{�1��|U��[�����$��A����
���Ї����AQ?|Z��JT���:��&��ئ�ƍ��	tE�u��b�)��!X�Co�r �џs.������=�a劫���3�޶m[.?�g�U�b��y~���勗`�`A��۳h�0�ƾ��I�$���?�V�B��z�C�vZ/�`�e�5�a�,�kHn����'�bsv?��q�G�����EJk ��)��
3���D8��:Q���~$~�#G���o����ɟL�f�����3/���bډG��`0��-i4�7v�޼y���ġ������7�ƂjR�z{�眳8޳s�o<��3�8b�fD%C��E͡+릨�n� ���;�@x���gq�&(��-𡹡�,�ec��G���K��\).U)�DīUث&��VQ%�P�����5���L)߁��*��&�:��<�D�@��%Ä�� �ے# u�f;�h@�)���UIʞR+AD*�Ry�?��n�o43�,g�ѲY�=��Y��%�R��BO<^�Ք�W�S땁��#��� �Uۏ`"+���9�ǅ��C�H������Q-��^��r��¼\�u�j��'�U��&%���ںp!��=�Q�+{Ԣ۠�oK5���Y���1{�t_*ۻ����AW8���ܱ2wvm����)�D���!E���g��t��	��'{�Zé��!��
�&lo�&�
�û]fyβE�0�u��c����X��BN��8@.wK��Ii2��iR�G,�Vߌv�t�nx�C��Djy��n��P�Ϯ!F��*4t��}�V�An!��-�Q�3
��d��$x
鋬|S=A�j�^ܱO�am�ņ�*�h�q��D
1/�M��Έ�&hm����,�Ժ���KX�5[�*
��`��״A�ߗÏҌ���}�l�:�}�a�X��C�_w��K&N��7�߻���.�b���SO��i��c'8�f͚n����c��j����6.i���/����x	KS��GU!@����y��mqO�}�&Sd����ŋBމ�+l�.�RM�AF���R�����h�������W�q�0gC/�8q"�+�� ����㘽/~�O1�����R�t�'���	&;vr��� �Wo�|��e{���ç癈�VܥJ��N��o��:)�e�P)l�*��O�y��Wo�<6�?}�#�.��{����1jOX(�~s�		�&FQ����שV�u/g[�o��p�?va.�4� P�3qFcKv��xq��Y�pU����	���{�)���@zh�s�ah��gr�4Y'���Ԥ���MI�od_q������/t�H�#�����ff�e|��"<����qM_G1_N�$T��#���Dxwj�a��N'b�>4ՀB���pC�/�0�H,�[Hn%�.:�S!�	Z�控�J�0\rE:���0V.V�,YR�=��޻jV���	� �y�[?��_�,����8h9����Q������{�vE�r&���W����J����]���d*"B�L�B5�>%��-~-<���WZ�ia�3h���i���#i�������І�۪a�V2��V+��������T1ig:���'�Mד�A�K�*K���l2��]�D�`/��Â��A,��!�d~CH���
uW�1�������_ ��,�����"��%QE�nE�hM}�9�v�+uU�lg	;�m�n��戚JB[吸�k��pm�Nj��z-K!QN�&�O���?t� ���ZxK���t�_=�1�*u��-W_�z����o}�[��X�z��o���@L���"��H��[xJ�Kd�-�:	���/\L�b�Ie9���s�	Z�/װ("������<���%{��A$��T�^\����4365�������Ë�DK-��׭����_]�n��B�\��ڵK��>�pwW�|�s(���#97Wܳ���c]��t���.ݸf�������\��Qz�@�\:���]��?��;��ŝ��=G^y�?��?T5+����k���O��jzbXKF�j!}CMeұDʟ��{�8�BaN(Uv ��R*�]]K����¤p$��|z>�l�����s�j!�̈́g���8��;d�K�)U
����5��[��QM��)��0�E�j��Jg�I�a���J)�QC)Q{T�x������t����!"p^�j�9?v�j}L��L��I��{�Z�BK�3b�\��o|J�1M#a$��i��K{0��L��ޞ��yv�H�zr�D�;�^���QAR�6�i�⑫��T����5��w3�$V�J��ѣFG� ;@Ŀ��+����b}�6]���7O�?�=L�PF��RK��W��§&���Ɖ�
K�d�"�q��%�mÆ�Rj�+ı�[DqA�˥h��v��m'��\�C :��2�EO5"�AUN�������)AĈ����S�;�F�H�RM�M�Zg�)�����]�3��^\o��wؙ�������V����V�I�kB�a����h]������o,}�>���x~B��ŋw/%�����C���KT'%�Ɲ��UA�%��yڻ�N�H����𲠭�ݭ�&LW��9wM�gI��V.��{�_+7�;ap�P|�r+?���ݻ�7O?y�y�A�c�r�7޸�^�r%r��7�����>|�%hy�|����p�x��ł�jK��"+���&G�h�&�'S�C�B�r�b�0|���*{���i��0р}MT e���oyqZ�U2�=��X�n��#E�?�:?��?X�z��4U����=��9�LOtI�{��9��߿n�yѢ�k��'&aP��j Zዧ�0u%��Z�A����ʔ2ټysO���}��'K�6lX��|㡓>� E�:;���.̚�!;M�\�WJ6$3!Hb��Ĥ�Or�q��w61�m�G����qO||bb����,�p�2��	���:55�g��M0�_|l{ix��[o�����LEw����.�Bs��}D'���֔�\�l��>���'O���������a�c7]L���U�T���5 L.E��=f��5RC��e�r�)#˲�7ntk5"(4S0�^޶��S�L��g��~������Sc����%%&��W�}�ݣ��0���;������G^ُ�S��V���
Z{��[��-���Ӓ��� ��z �6�
I0��\���%LS2	��'�5O�\�
�DS��ZD�W.�v�P��¼-�?eA��?���<��wp;ZgE���I�R+n܌�
k��@i�f��Z��o���T"u%(�!�?J�j��KJ�Fq0ߢn�jif�+��ގez�QLD64�����p,[t�·��?H��@j8��%��EX�=B"7P�3�ռx�0l#�I�R ɥ�������߈hA�^��;C��L���g �bQ
A�\{O�+7�{j��4�pz�,�+s�9L¡�/����{ժ���_��C�&�Ո_w���[�=z�f�a���~�������e�	g�]
<�!���	$��EN�g�m[������a�.��cW+-���,-����dl��3[�k��3��L�J���'�}G�k�����z�:o�Z�a���z���#o=�L�;2qYU.����|h|jj��s�U+"L-����t�����ر#_̻����ж�]S�D1k+dbT�!!1yt��qɥ���L<ݱ��_<<1=��ґ�Ċ��v��}x�7G���ٓ]���n9����*C�s��ٕҩU7U�G��HhF2��#L�<gt �!<�A&�v]|��8�8�ұ���-@,p�AD+�U����N�8���@�d4��+�ZԦ��?9�"�|­DjsY�:����職�<*%*���p@4�e��j���5n�is�L\y኿��_G����Å����6$�q�!	��{Wܴ�"��=�a6^p>�֑��)q�'; Eť�ƣ��_�����W��G��J���߶{��u��b���5M񎌝x�=��Ki�:��7�B��޽�d���~���ggg�\v�S��T�������\��P��9}Z��9���
��J��E��AM�S$23A�����F[���Rs�����x��b�#�݆$S�F�d�C4x	�+}\f'<-�o��$��Z��2�M�2)?äc�Ɋ/D�H�Z~�0~�g�c�
%PFS����/�]䶢�0B�yR�p�_���S�aj��
�mQ�Ul1�e�{�&��*V�VD$�.SE��ӧ�Y�дB�f��i#H������&�1��6n��d��Fe��G��Њ<�p~���_
�\.��M� T��(�����U� c��	`���q #3�f�J�J-F5��1]�0f��i`�bk�r�eCCC��v�m��7v/_��� �n���E��(^��K/�D�]��1���t�����]�%K�N�#�j��eFI���e(	FrhH|v��F�W@��P��8�4��
m)έfG-��0�����&�5�˘7�J����u��m��w1��:?�я0@N� 좩'N��馛8����.z���#�<R{�5���I<��-���1>%u�������c`��!s��]�)b��(Mvl�r���7`8�p�O�o��Q�B�g*N��h�"�˘[��\�����_Q�d5(�W���,o�w?�#~�U�p�U����Z�nO��eN!A��6u�ْ�E,��.�K��1�.���?{/7?����W_}u�"h�������������Q���<�&� f��L�r�����L�}�����w`` �c$�}$7iS��������8%���U�VUk֯~�+E���U�^� ��M�Mձű2^{��|�p�]����c�/}�K����&�ۋ�߰�<X���Ķ���ǑIw�{g��M
νwЩiٿC�S�z�͙N�q�{Ţ�"]m�>�pD�j	���1Z��r��4�`�=�P8Z���F����Uߢ*�u�B���f�O�^�o05�p ⨾��e�
�}�Z9x	��0!�:�t�
��vhK��l��Ia{��Z�át`%�SLͳċ�.]���dJU��_"�nҩ��v�"&��2#��]R4Etr�<��En���B1L��t�����t��MMMFMɱt��Md׍`�0F1d�`j&�WԦ�" �PL�5��FU(7�Iutå���'� ��Gpzjre_�j�����e�2��'+�3�x�ꥪ�l�����#��-����9��-��w�������_?�r���.<�o`p��}߹��̘���lW���-~�(!!1Y��[�q���d�Ά0�T�1�d��|`� v����B���1�k�@�O�j%l�����@(wuu�ċ�a�Y��}E�aMƁ�F��↉5dؿo�׾�����/�X����_�k�I8\t$(�l�Z`-[�'�&rj26S��;z"
�幆�rd�ڰ�L��A	j'3J5�r�R�2"k6����<���'Y��?95c��un�*T���c�d�\U3Ij�SI�@_/�5�ޯQ����("��ӨP��j5b�����x�tl�R-<ǪW}�1Sm�e���.A�%�:V�Ϭ��Ч\Ѩa�Z�5�8����T�#C3tY�#Q��ϗ�g�zAq�T�Cev�b���!d�S��Uծz���K6<�f97�ח��8~|�ꫯ�T��W�讔
�J*e�,����ꁬ'��������3�#th����߽���d,m�S�\WG��_�-#������^�R:a�m5����l�_ҟ�������-�O�������B2(ib�tLH�����L�K��\�����o��v'�dmgT������=�rY��?������.9~�^7c��fL�&���*�6�(A�Rnw "�T�F}7��a?4dۦ��j��3U��d_�@)S��T��<U���i�j���F6w][�>=�o��V�g��7J�RG^#��G,��tG� k`7`P��g��	�X(G�nh�yCϾ�j1�v}(�Y=�����;����oC���F��_�۱��1�/�'74�V��0�D�Jcff����f&OQA��bJQ�<��-�kp]i"��N�j�"�j�_]���(
��Lr��3��A��.��$_(��ggE k�Ɓ9'E�Ծ�^���9�p�8P!�k���WA�^S���c�=�p�֛ #�؇��[^~�e*�����2/�����0|n�淥`�12FU�9��*pQL$�帜�Ї8ۇm)U�yJ���x���"R!���tu�cy��~�<�Դ ��k֬��Q\���.wn�[,�j���MS/K�Ȣ�hgOfO���|��.ޯ7HE�177w�歟�ԧ�}�!�ۋ/�HL��]�����^�P���0'��M��zUb��\����d�{�<M���9�jUzc�6L�֫��C���+��[a�����{���ƈmQ#��[)0�.όh�hq��lW�mT�����!�k�g�7U�c�76S�F���iv�n&ss�4�0V���j5�|��W0?,�����n0=aw"XŅU��x��K.��z�71:|כ�L#p��ꪾ���k���?~�(�0����S�O`K��p����e�M�u��-[��_��L����\չ{rF�D0�b)�T�LI�dQ�β���g{���a�g��Wk�y�'Y���Z�l��DQ�H�b3	90��sw��j
�x�]�ߨѡ�_����ߣX7fIaWt�3�/`��^^����`W'����p�
�lnn�?��M{n�^�����鴬��h+aۢ�Ià#zD��+	"������YE�@�oNF÷T\�鲛���b�W � �/%D��pwX���`�M�Fy����Ps���u���I��/UKX5M�E+�_C�B���(�*�'߶wew*)��f�k�1����W���%�����	!b�u̦+�v�������JDF�	��#AN~'�
��&rXU�D�y�R%�N,(&�	�7ϴ+n1�I������OӂiJ�ҀO�ʢ�D"��Hi�#i5~G�UlC��#kc�V�]Y\b	�Tt�R�u�!���b�)��9�_GT��7��{�פ���~��n��S/Nϖ��NLz�n�������˿�$w_Z�������;�� ��g�e���ă���)'0M��ib���00=0�����!��d8w��x9��}L������;�IA��9ō$j@�p*���R��ȅwE��a�Xk[J.�!�d?pͦ�k�F�~���w&�`����fwg���/�RX^w�ر�c��α�����~� ��9K�\�^Z�&T;�6e]G��� =�%�$e%p�P���Ϫ��Cxvz�,/�{�3���������,�� ,�|[D0��V�D!G*�3�:;�;;�֩� � 
��ٜbO�L-#90���9��j��Ѽ�r<W�Z)ה��*�A�!l�Y�.�[IN�����Yt�9����j�S�aZ6|-�k�e�X�¿�w%�>��[�ή����{6dó���@W��еf�d��������	q=g��͆T/�k�z��o p]3<_�R�X��H�T�Ҵa�F:ea�-�~�j�v�͋ss�Z-��Vd̗J�ꥲ�uM#Y$WƼ��F�Q��/t-���ơ�S�+�&�+р��[���h�ũ�)-�g�Z-���(���i����Rd�	S+�G�LQ�x-x��(6:!;R�2k��i�;�2 ��JN��̰D4"��.�Kud�zjRQ|��P"��5�}Gq,#p;���������TAv�/�ʮ�0S�����4=�k�i4���ܕ�*� C���haO����N1̢�'�(�*���jq���Ith#��k��I@>��@��0�YR���(a�	0v o\;t���s�������޻&�_}�}��$�~�cl�i"_'�$�>(�<�2:�7��!X�P�q����ETqr��
��۷Rց�*P6��j�^TG*�=�4��

�3#��]�p�7�@~>Q������k��ܹű��>�,����AV[��H�aI6Kj&��b(N�$��^�+@=0K�Uv!�5�a&2������.ov�D��H)� ���`]8�[��QVL�:��'A�s�����"����B�� ��Gd&6��.�raq���o��/��\(���p��w�l4����C�� �QU���:�e����k��y�A c	%��]��������=�K�~}�s���Lw�\B�_�[����&�I*͵��򩲌M4ސ,���������ӑj��3��׋΢������r�&����0�D%�ˣga�m�����k{�1�y���[f��!�U��`KN�0�g�}v��u�_=�_�]��MK�=�I�����_� ���J��. �];w��JȘr_D����PJ`#��'�b���A�_z�%�"��{�����U��zꧻn��;n>�b~�;�q����,1�3.ƪy�8CQl�eRG�M�곆'�G[�M���d��ᡡ�\F�S���I��ęݻw�S�d�
|�W��Hs �h���9rO\��~� |e��m(B����'�9�<s^�X3�.Maմ����a�Ad��w��W�(���snt����,�%C$(ݐ�S
I�y/F���i|����$�|2����)�3�9��0q`ȶ;s؉9���ȶ���ݩt����1�54X�`0,�.M��#�
oMG4�E��
����_�n��V����؎m��r��jW2�\L��$S�DH,�K���` d`
��
��M����]z�'�A���M_�R=_��O������7���[��o<��G/_�T�4�Ҙ>RGhB\UG"��7q�ָ�/(�C���*$�ôNl0����-�yvp�p�@�^AM9vܮ����S�'&>x�i�&Pl�u(`(��RX/-~XIN۵�բ\�  �e�����pT|W4f>�ը��F>��3I��ɳH`������j��}ex�.	jx��_�8��� ��x��c-(.�$|�"��j����������3-�V.\����D�b	 
AOW���L�\ƦN4;�$v�sq4��M�]	�B{��K��x�zf�pH �U��}ޙWI���/p�"�\��nCIa6D�֌Bq9�=Ռ�� ��#пi���p��e���m�?����s�7�tS{[~��wj~�ӟ��p�ܹD����|Oo�
��ٿ�p�s��0��J]��&Lwn��~b����?�3�!�=���vJդΒ�K���@Bc:�	#\Z);R��������w�ygx��tw2ӝNwMN���I�gj":ړ��h./*z�l{�,��\9�&k�]����/j���ֳ?����Y��۟���u��ī��5��#B_���^t��l��]S�n�%�Pb)���zy�P/wd�;�J�<3ޕHܰ}-l�C�Xcd"����#��݅ds�����-ݷ�-��[�.d��V@�hh���U�J�`=)�≷�w��k�k^�m��@&��v�j��ۆ&o���;�a~Vf����T�0����/qQ��9�&�R�!�|�f��b�/)������_@�+|����,1,�"1��$����aPTNh�M���0,Ȕ����
$0ԕ[�a��|�x�*BXp��ب���[=4E-�i�U>a�&��b����jd1�?���Xz�H$�[0f����2P1�zƕ|���T�n�5�nݺn]����Jݲ6n�?
���e��m�8!n��/��ȽN�Ur8f�u|���	�un��>k5��Q�n3�����{V,¤�K .�4J������d�
\�`��Ǒ	�8�e�Ǉ��T�0��@�l?q�(��ф���>���ONN�嶞�̙3�ON����������`���;�P�~�mI�y��`K��,��yK`qj�2A]�
�p�����Y�{@M��
l�p�"�ѩ�;��?]-�<��EԐ�_S�Pk��!$e������&1/�|)�%уg�}��E�~��������~�,��`м��+�Zubb�^��7�~�:�d�~[�l).-OMM�1+��{�����7�^���~[Ӟ���˿��0�͛7�<y���9��al�%��fU3�����9�$	��$�E]3��22;	���i �TGz�,�7���a{ù����w��|��sO>�$�`�[o�|���{����pَ�AJY�e���ɵU�aA��5��cq Ȭn����H��@G���R��}��@|���n��׿θ޶�r�U/�t&h(��c�x����텡��֯��w���wW�+p��l�J�ٳ��g��.M���*�d7?���A$���\���?�Q���=oY�E3=~a~7KN�* �ET�,w"Q��˵!In������˙��p��yl'!-�|łe�Cd01./	2ǻ����5UU���6@v�R^��Z ���KrM�Nx�D���(�/�:�^0R~ݜ��D� ��UWlO��..,��4|Fsz6�J�td���Q��z�q���k:�<s���?������i�zB�0v���?�rQ�@���W��u;�C�%�)��v�X�ܪ�Bz^�1�q�4�$�:� s5�����+,�H$�T�&�=�.p�+�����Qc�|5�}}`��	g"�@�mڨ�&���\$:��.�%���z6�]������W��+_��{�:�����{�o���h*���ކ5���u�j�Es���ӗ��x��L2����j��2%C�ڰ�.{EΏ]�8>Qm6�T꩟<3vq��W_�]�-J���"2�X\�0������_�L*	��M�z���sEJ-C���ݠ�#2}��X�p�g\��jK[�#D�(`�&���������UT0���T��P�rS[���~�������9	i �K���K+�Ξ�ŕB{gt�����+͹�Bggϥ�Ӫr|ݺ5s˗.N^ݞm�vJ���6�Pg{���N�8822��[�`>��!o�}6IgG��%�@6��$L��]�d���tk�����7�9�](���v�ȹb�?0�L�T'���+I9U0%	C4���%��Ͽ�V�����|M�~���w�����,����G�xvt��FR(d|G��53N�Ÿ���	7(AV��R�C`��.l��Ύ�L�2q^n�oڱ�÷ܴ����d���=�I���b���'FGGO��S��_����ѹ���ן8qB�m�c�-�}�Ԫ(djW�Y\�.�l���g~�;)���ڍ[�a}�p�֋㳯����k��v# ����;���rݤr�8l�0�@Y�Ε��mKZ��x�i��cb	,~ȱ��� �`��r��0�~��Z�0� �e_'�]����ry��W�T��H6` K�a`ч-��4�е���_x-j
�D��t(Δ�l �W�[�ȉ�*����5:� .Y���qJB9	�}K%DF��y��H��� �,TCMUT���1���܉�_~.�K�]&��˿ ��ӳ���4;�L�;A��y�>@N�efX���\]�<�B��z0��ѠNC裇rj|����J�	: �s��1)W�bs��Ef`�?kn�nf~7�K��6��"h�u��q%Z�*��F6�!X�Pڂ��D�z6ب� >"�%P��=~�+_����O8���_䨥���)�*6��w``aa��ALrQ�s9�U��J����0g����SO��?��0���o�����¯�v������r��2���Ycx�ṴK?$�je?���j8�2������p�#n[GO"?~���k�r�S��sx}�g/_��� !�\�t	f	6�ٳgm7 �ښC��k׮�=`�>��Պ�U�x�	j���#�����ؖ#���q�?~�.{Ml�*��,l�:U/�jXY-x|��p��E��rEr<e"��x*���+e����o0�O�`5ϝ;'�.��}�{��V�5��{y�G�g�� c#�&i6��>"�$��-������΀��x�`�'���#O�r-ꭐ0����M)��>|�0��m۶�\�HvU��	b�pxK���.]���w�-��[�&�0�F����];��w���ep���"���Z�t �˔�s���#}��Fj�m|����1�QE	����"�I�"�d����à6֑�].sn,O�n2y �d<�T��$U�����7�R�� �P����l ��9	C+twê��A�؂g5��z�R��i�nD�*�(�R%�N��P��B���W�w��=��Du�/z���F��j�+���L<�"���mzeIU����u1�$������:7�cwogRQ������Ĕ��:r^T�Q�8~~��#���F"��z�	���ݕKX���9
�kXJ("?�c�&��]�x>�aÆ2�'��j^沆�199	��!�8���q���gqj�2»cp@�Tt,�����.�E� �5�� �:}��Ϸ��I�]VGBrm2�%'��ݩH���Hx�aMd0�E%頵���v�Y����dG��J���G��άif-7ӻ���d���G�v�����u�.��C'�8��P�K��R��	EqɮWW�5�uҺ*$���swa�_��;;��~��������wW*)�\�3�<��[G�J�d��KjZ`hR.��5�`z{{��yY]�F��H�߃�Z7�I)	҉d!�3�R�X�r���-�@�����cSIl�f.�ny~ ��\!�N��t:iY�|��s ����
�ܖͺ�؄YAU��d,v�0�K3Ei������c�fI�i�l#�%�y�����)�vOҦʶ�'������+r*��pU��L�Z��iz~�$ҽ^*�^D[!�`��&F�`2�J%k�V�f�` ��YS�m,����ӕT��&����T �w�*f%8uW6[��XD�OK�Ku���#�f`��1J��R��d��		w��!�����P%"F&�DhU��e�@���R��@��P�0��d���޶���x��k���/���؃I4���G�a�9}�3C�B��-_�Ԟ��ѓ�c05��I��i�zN+/,i��כ:��S�i}��@(�B�5T.Y��cu&p<r��S�-����i�������^�Vs]�ᬭ�e]�g���V��r˓è!䣯��G��t _<��"�2J9�]
�D��;!
@1fa`�@�(ulr ��v;�P�����+5������^�#�3��J��_9�b�[	N���\�;?F�bRȞ��Րc�ˏ,'�>�cҵ>9@���$��;˲��Z�svv�+�61L���Ԉ@�XV�����w`�oa�7�&_c5c0��q���U��Z;��������%>K�� �ͺ�å�^�n�ǕN��^�����mR \aiŧ]X}kuE��9_��P��R<]��"��497y���J��nYYYz��&& �i�Q:��L�F
� ��!FFj���{�n��1?o?��C ��o�hn�cp�}���ʁS��mʣ[|',���tq�p����`>w,8�=P��i�EI]M�~σ���5�R�e�}����5aK�B�1���KM���B^�b��-Bd�) {.|�V�ժ�V_Ƶcb(ld�N�r��#єVe�$>��<<�ŁDb�J��FW%�� Y}@ͻԙ.�P���Yڰ�p挩hK�$� HD��e�t�|�j�Jd@��>�BQw9�֡>�`�c�Ʊ�I��ٵ��$�9<<���yr��;w.��g�������_[;���������hY9y���������T#0��w�}��_��_۵k��g���W��L*��:@[�w��o+�ĵ5[�nM$��,)2�C����ws=�'��Eq,�m�h��q��AX-��,��)y�c�qV�⏳�!��r�P]_��g\�����m 1�����mdd��͛7?�)Ȇ�SHVD�#�j���J, l�ʑ��~4{�\%�ᑋ��1�����?$j��6��H�S�gM��Ua�3�t"rvj�2 �N .�DR�=�=x��,�W\t�d3)*�Go���,��Hr�U��/��ñd�0��V�G��a��{mmܜZ��+������ ���-1����%�����,����z��[tP�H�\F��$0�ʚG��VW��y����iR+��3�j�	��Е����T,.{2����K��#`ǔ���z���٠諨<o�u�$	CO�N;D	<�h{n��l��{�������n��s���������o���_������7�C0W������K"@{ ��Zf8�}��2�Z�	W�"�[�+\>�{���d?�^�8r1�j� gAq��yu�_<kzBP���T�Y9�.G[�*�B�~�%,t���aY�(�+�GX�#����I�bQ��d����i��RQ$˔>Z�h}�DDA ̴]��Ч�9�0-���PJ���9j��U%�V�PbEbKܶ-#*�Xit��@�l�!("��E�4A>M��I.a�8f@}*Բ=�"3��j���� �˪
�A=b��V+�����{qieso_{wO"�Mw�^`KT�\,��4LҒU�詄����m۱����'���}5��$��Ki�����`�lܲ�|f��IlE��`�������p%�j���~n�r��沘��(:]�_�b�A��̣�*����|q1-��oB�ŋ�"��a~�?�!�#^�M�?S'��"���f^P�P[�V�i������:�_�}o\�x��=NJ�����AKWQZ�Jy./'�DWYQ���Ub4�p�X���0(˾5á��B��(�l��a���Lj��������aP(��L<�� [G���+��c�E��b�'D��gM`P�k�[0Bx.�G^
��
a���@�/�?�%��7�*�(T�����H��C����.�7���G���/xO�Wd���[q,�}z]Igg&�@�mlX����T�:L01(�AtóO��Z�ᶦ�533C�Rd��;��I��� �A>������WGmj��ԡ�<Ν����թ��ǵ�~H�y���m�B6�����*�"��E� �3%�xeY~��ض�ہ�U+���P~zSո"D����b�3ޚ��7a�]�H��pH
�z!dl�BAو"a�&U�"����))s?.'��A�K7�)d�
�:.���T�T��․
�f�����8��6��r퀀�u�f,R���� ��ߏѸ�7��î����w�V�0J�ǽu��6�_�S��	�Z\g���a����mڴ	�[�o�����B� 	r�``�&��0l��nl�}���\� 0���Ijz�^*�� �󪑋&"]�F|��.�L,!���l�+�
|��*oeMŝ^��.��p����R�І���(�-����X3d:vw7�2���|�׆��R#`�˚'��(�ԈC�ٚ[����U)���㇢���A)F�s~C���S��@� L�L�	��+�Q������GP\Gr,T���@�����ߕY�õ<�;D"�%`40/$�bp�\�\��l�����H Űa0����o��X���_!I�E2K�8�t=���A�Ĳ^?H6�].�F�i�M��k�T�l`�H��Z�U\"1����>>��)�z���ג;�wa}7��VVj������|�ɜ���F���NT�����C^Y�1\ӳX��*�۷���|�\�t��;���tu������#���'>��W��4&V��=�銁���><d����QD���*�j��1B��}�@�΋R阒$1�H ��Yd2g'��b��T��kV|��Z6�#�f�>�X��3Lp=P�Aqy����rq� ���$�k�K�N�AnC�������(��K`���L �X��|�)W�U	I��w�e�Ĕ3��M+cT������
�w��J
�0'H�)���F����S���Ҫ+�U;iP��˦�&@e�	;Ȋ��۴`7�QTl��RsU0_��}-�fC/��'�7�y[�/��&�w�:5��ha�7����k���+�z�5^�2s�|�'�8�7� �PTg�*�}fn�/+ɆҴ+�&�WeIC����8.�i ��r�u�	D�V��kT�uծ�BP/d���`%$�>-1��H����H�GL�:ꮒ6�0;�{�_�W[[��Re||�H��^�AHMLL\�t	�|&��E��ȎiQ�Z�arF-^�sx�oPn\2��]
�=�c��|����݌��a-��~,6A-�5����;�Y���r�!D�[ELh�y�$��mUd�8�.?"qA��������I�O�%T�h��g�5�`E1O�8{�}}�$��CV-�G@��>솄K"��� ��ݾ8��3G�[x@�B� ���GA��}�v��u���P�U��?�8r�D���T���d�7�V%JA�&;��\����0�\�8Ǿ}�������x����i������Z����_�"8d	%�q'Ə�"j~��*��::���BL;Wj�������Ҳq��3��^!g;u��[\�awW�^_K��1#�5R� V�}%��`i�m띝�dC5��C��g��&�G}�N�r�J7p
�Lez���a��[��2����^X�E�Đ�� �AK�u!�i
K�|V������gvx��ă��!���$v쐱t	j�L���&�df4�+4ke��U�@Ϲ�a���;w��s��=�����:G���r�a����@
�n�X�|�ؚ�<�d�j��l��`ki�5;;�c�晙1aEt�
�O��a�\�ev�sY�2qr$�g(�W�CXD��ô</�Qƕ�Uv�te�����������0�\o��B&}yzf���s)43�B$�N9�	�JղP~��v��� yRHRg!C���i�q��*��Vo�tr��W�M;*k�����ߺ�R	�)TM�H���R�$e�u�Aj�
�#��t��:>����VXՒ{LD��/���yQ"�/h䈋�%x��ɉ�Mz��a�]P����^���F����t�Qb҈�L����j��B�>��@s�w��E��|�e���W��ֻ����%���mܒhHV/�4�K�ڻ��Jd��<����RJ�zQ��*��ͥ���ɸ�T"�Mr�Y�~0�\��&P����}�n��[�7L�\z�����,KS˵�~��p���<ձT\ɴ#a���Ff�v�в����7P��MS
)O"�)�W�ycG�%V���G��eֵ ڈ�Fb�:������N�\�7�f9�]�8������D 4%�g��Hi�����0!XT%a��cQ����� �=ɀ�LcpX1*��p�D@��3+>�x2-�J�!��Q����-C�-0Yh�@b�%��H�#�ӡ���Qe,��+v�6�)oq�լ�fR������@�;�����eEj/.$(	ĭ�q�O��{a�ܶ���G�L�K���\)�i��y�us����twz��N�P/��TG/M͎�.�[��jy�/���y_��:4mSV�m�S�Ҷ�����ɺ�g:���.\����̪���_9FbHpUMxM���ӂb�^x�`�r2�v9���-n51�ڍv�g8[-G��:�;���fG��(^�H����Y�?"�@���B��PX��a��_d[�&����###0Z@^��g',�9�m��033$��� �DAl�Z���(K"m|RK�5b��}%������Hi�~,����(�-��_���3��IC^ᎃ [qR|�h2��׋2&uLl/�0�"S1������O��e��B��
�� R���8gsa+I�dg� L�����+sss���b$'�=_9�N��Jnօ�F�Շ��#/H=,s�,C���&���u�۵W
A����x��I\ږ[׌������}H�A�gv^�M��iI:�
ՖF0aQԔ�L/��<���?��#o�{
S�|<#9#���/��ӧO'�9FQ܃����l�:^&D
�&����aG�8��mZ>>��0 ++x��BE�z���5�RS�ƽ�Kv`@3�m#=e���qi4�T�u�>�T����V�PGOw/|��$�C�rt�x���x�&
e��5�� ��N�}^St�CSp؋�*��S;�p�3�����h!ӃΌ�������l��a��n�˯/�&���?z��|��<�m������h�s���;
l����=��q��t2�K&
�Ņ�3g�4c ��`KW��a�V`�u��|rK;��j`R�L �,�>�l K@���ҥK�������J�k#K���p9���̈�㣰4l�1�ʺ�}�e�L)!#��~at�ȑ#6l a��~N���]v�FH� �	�D�*/���C�j
fR	���V`��{�� �X�
����+���D<G�sC� )ַ��!G�N���Q&} �����G?�qp�y��KHUj�;��m�d$K�VG��j��O�-82�>�x�]L��穪��G��/��d&�Ȑ)��*�\��h�ۚ@=x\2��E���D6��������e��oy\1m+�J65�~>�t�i*�Эf�\]�� ��;n�a<���p��aQ5�����RL�"z!u�H�|~����TKԶ��Y`naV��	>�*7�(�f��Nu����a�a/��2� <��r__���$�!���Ԭ @�QT�i�"LHWW��&x{Df��u�T傋��Z�:��5��Jj(+2��j����`���0����_��s������@�-�M.�����|�L2��PZ�l%�*��=m[��ɋ$ �" H������C����s:��ڵ�\AuX4Q���<��T��]X*��+C$e�\56��+���xt"��
�9���� �oD���/���<����k)��A6�]��妐��S]�z�i�r��8�@$����ߞ�|ۍ��;�5����'O��;0ԏ�`6�3�+)����
���u�ڵkA�==u֞�(���g����ߺ��R.��K�B{a�a�rWˠ$��ڷo��_\YY�"/S*mںMM�w���> f��!�3�3�����5`Z���S�P	L�t8*�������M�=�f�����p���ç���>�������,�E��?��͛�N�����I��v����?��K2�]H�aG��냃���ҏ~����8��$rC��Q�4�5z�W*0�/}뻏~���@�ى�J*�����i��'���\�^u���''&���[�"$���U�^���٠Y+-,lZ�3����df�RW�D׺��>v��K]G6�H���h�:5_|��#��F���]��?=79�p�nae����|>�X`�i~�Ȕ��������{�l36�!-�;�Q)�Q����Hy��i�\[=�8��JBV@[��d�!<��S\Z�1Ԗ��;{�^�8;==�$�9d����j
�@�ڼ0���������z���*�ݩ�Q��[Qt��H�(���ٖ�s��r/8p��G6mz�����-������́<kk,S	�!��_8l�,s�X�U@)1ܷ�Sz@6�`��Ϧ!��+QP.UMHz��qA��/R�5w���V�%���h�D���U������0o�J{�%���T�~�l�K_����o�s=���� n�
�%_Y\\��IfU��]�@�g���.�j6 �]��[�to��=7���j 8��=p��*"��lX�8����|l^{�0�bU8����V|�V�j�+�"��*<�L=6�#+0ʕ�\�Q�!���|D�D�ϡ����t���K/���=}����� �����0�;���k���>��'�m����E(|�ܹs>� ~�󟇥y��'�j�������0o��j�f��h:�%�X�J�n1.���#� ���
`���G����ˇ��a/�h�G28ES�;/XVP.�@imܺ>�|��	w�q�KϿp��Rz� �q����+ȍ����w��ZzO s��������|@kVd�i�2��]��"��o}�[������!;�byӦMm9�q-ת���s��A���N|��_?q�4̃/'����J��`�ǅ𭁮Ƚ]�^IJ��~��;v(�76���܅������k�y�e�5��Oܫh.�1��K|fx � dD�����!eq��b2]�Gqg��2�H��[$+c��GO���
�G�j��D��Z�3�5� "��z֮[W��Iq��(�0}LDIU �;��`�Kj	 �LNN��nI�c��U��1��谧v�"����n+���+z�|q��:v��}M��ϝ쉆$4�@�]�J��<�w�iav�[�54�7޾{�F�X���n����تb���hZ,�#�%Ƨ��,���Y#ϾM]}��b��c��2��O��F��n�3�a�Y�5��J��l�� ���m�
����N׉�R.?z��EuK1���{�[%��?E��p������|��76nߴ��_{����a�����s�C��r��HF�,�*�N��k6Z`^ h҂�"�>BI�N�Aa�L{~98|�g�}������J�������{/�y�
ם����c')�A�<��G�Y��Jμb�!tFK����;�I�H��I[�.:b���E?ܒ���le�K�(k�d��a-t��B>!$$�c�ݫ/nh���={����g6|�#Gp�f/W볂��(�dJ�]��J�cg�>}z��>�ɕ���B�Tr������&*cH�g�k���.�T=�&=�kz�	B%��󁺴4�3t��(	�5CmZ����w�E�6ߴn�P�ёR��Bi�rW.m7�t�1W.�._�I;^x��������#�./�7���!�6��k�c����r7�=zt�?�.�/X�3#7�����{�W,�ٻw���oZ����~y�'�J�M8z"�Wtj�{Mt��K{׈ɶg_;Xr�/~ꃎ�?t���	��G�%u��w������|��7ul����
�{ߪ�uU��Z��kdx��ĉ��5)i���*�ڙ��o����n?}fl���#=�ֽ��Z�����wٔ\%��s�j�'	�i�_y]�`Zԍ��F�BCsՃ�d�`�UB�*m!���_�=��B��W�}t�Q���sxxl�W^~	�>�!(��&{�D/�kv�K����c?-��]cA�k��?{\uJ������>�Q���M
iZ��, �zQ�s��4�]XXHi������������;��b|2�����J�+�h��;���׹����fB.�b�x`؍(�y3�L/`|ĩęjq ��XӸD%/J��qqc1
�D� �-�%��#IJr�;��������~���}�s�Jm�֭��6�'�/|��ѣ�QCH_�tr���F�Q�	��H�>�Å[��/^��ꫯ^�Ώ|����9��o{p��t��g0��@wxGDT�I��F־Q/39���NCz���vr$�9z��o�Mk�{!�%�HQ�^�B|���;�����t�����dR��N�����ٳgo��f���B���[��X�["e��l�����@�\���6k�����+�2��}"�����V���.XO>��'��M��o��xhl�N�ʶ,���p�����o�U��8qb�}��=��� �A\�����w3|fb���.�����[��{��1����ڵ~��w΁���FÉ�`�j���YR�Љ�&��?~�ώ���{o�v-\?��1RR.Z}�ߎ<xp�r�����ǉ��+e�S�R5 ����&|���R�V��|�=��J�E!�
0*����ssE
�u!e��ꗎ"T� x�c��v���(Gig�T�HD9$�A�l$��#��
���8z�����ߴq�<��������y?�>%Hyn{g��Mh�d�2us�D�й�bf<��"Q���Hl�TH�
6	ʋ$����V
\.�I�)��U��!k�a�'5�T��WϠ�M����LXvR�3�A �82ϔ�g���ܔ�4�,v���ۿ��#���!��
�iK�tR���{B��#Q˹��'��a;�n8U��8�(�����Y�I�k:1ǁ�t@�e2i
�&�X.�%��Ex���o@��!��L{�冉�	���w]QMK�$��ĮDJ�VÚm����O}�S�w�3��'Wfgg.��cy���w���-w�;7�L�[f����*���e�@I� ��F��W�ljBԭ���w���`��g+���RݲW*��	Qэ�e����l3��-P��)�`�ql��Y��o�j��j���P�]-�����d<����v~�I�^Q�B��+P#0��t���,t����A2�U\�^���h/�?w���#����gOn�
{ziy�AR�L.3�7���_�,(��{KOg�tǥ�sm}p��6��-�,+�B�4�0��n��:�F�V�ff/_�p&��C���R�
��es��������yӶ��R��e�T��43�k3����t%��B��b�Ώ��G?�+0�+��p���=�ܛ�6o��[6nٵ}��t鍷o�fǮ=�/�کs�3�T{�����{���b��|����#�: )vCWS��W�hm'r�+ML�,c/{�{�d�+��������j�}W@L��u���۶����.#c�m4��Y�^����M�N<��^W�P&��H�n�~�#Wr�=�joɸ��4::*Q��2�Bx�o�6����A�r`�&T���Ť�"�����������WRo
1�(�m^�0��*��� L+���UΟ�Vf@$��0,bD�����p�̙3����빧�.iEz��7SV-�^&3��m&��(%n���rF�c��+�)ȫ�Z�g�sίC�aVѪf�W�l�� ��ԾP���vh護޺��[ð���?���AV�kHCO_R��|Ax�4x�J�K� ���(�+��5�JO�����ɂ>�1W�s���ú���<d^H��4��pA/\3���s��o����I/B���p�����9>� �y�d�m�����|���=0�[6�0u�
�k��s����>��u�]wj��3C[��k��͉��h�:���a`�YQA��݉�
SՖ*E�azDKފ����c����t)�׏K��I4!�N����bB/WS�V{�Pވ%"s��"�b~QR�5w'=��O��}�v.��(O���z�ێ��d�q//�J}���C�$���[�l�p��Ԓނ���Ĕ�j���%�_��ultwu��g�z�fMӋp:��^TW�f�QV��S8Ac�Xb�fO�:���~������g>�p��������[o�Y��U*#GD��nmdd{>���Ω��~�q���e�*ZB�$<�B�V��nOjL�{o�;q�С�S�9�P+O�Ncx��Fؠ��l��zF��ΰ;�:ྸ�;��f�ddd.;71{����P�.�D5u����XRN��&�d�zC�*kEeV��b�#�f�6���b�rȱ%����X���R�A��<�a�(����BTB�N�2��_��'fq$v�|䥁�/�ps0���^X�\W?y�� �M��ʢ깎��Kf{P ��7�i����#�3�'Q��ȘL`��W/~�\X|��\�M�ld��ȅ�(��Z]��������}�%��<��cG�w����_�?�Q���n��d(pP]4�=�}>�߸V�r��PG�LX����aSuN�@�CX����ǲL�"AVl0�7�b�^�(
�b#�Ε_�U~�Љ��
dZ��o9���K�bw�֭k֬�X^F���������������?^����woٺa�PS���ӧ����알�qb +����!���(�1=OD�PAId򙂠�������B�٨Ԫ0��-�w3���ROH˛�4=�_��Xc0�ᰰsc��#��\��F+��U&�z�r�U��~�˂��a����-�����B*��RZ*W%=�\�_�?xi|��R�� �gq�8��u �k�4;����;���[/�ZM�����%���k�m�fN��侽����r�R����������Ӳ~�wM'#fz:{�S؋�hU�&Z��lRh���y�ӟ��Dz���3M%��$S�rY6rJBl.W-%��K��;��ۿ>*��`�4�.4U����]�YO��:��>��R]�)��5AI��J�t�Y�TK������鮻���gu�u7��uh��%����+��h�����P�)�M��oؙ6͒5ۥ��*`�	F�;�˝��'j
��b�ؕ��LM��N�r�ԉ5=�g$	]ܼu;(��sSSS9��0�t�)�\����hK�@q��l&��Y݂#)���	wFD#�I���ՕɒI�ȫ�[6�x�\�ؗ�GOxCaƧteW�a�c����)��d���811c��ǁ3ȾЊ�k�+�F�Ԍ�r*`?MB[	����������q�kKѴ��]��(�D����Q!�;���3�����L���~�'g�Xܻw/H��~zzz��9�.^[����'~����3��n*���c�
��@�l� ���.v	��P�@���#�X�Q�0)G/�un;����!�S��ܹsjz�*%�3�������6"�(1�JEy�iv�����r�-w�}���p}%�����ۼ������]2%4����?���~��S6qCbD�����A&" +aT�t�}��q�J�a�^|�E��W_�+������	C���6�|��̲�����T �� �T�Wf���Q�+�(���s��޻������,_��Q
��%����Ӣ����DRgGj~~n^�� �y�5�|�k_{��v��z�}�}�O �\&�j�O�^�w=z��G��,--�U��5Y.1��׮]�C���)O�"G�o	�ą�p����6z�*�Ɠ��$�A-,L���5d�i��ђ�Um`5�-�5��6|��ѣ��]��Q*�� ���7ޘ�a&���$qL����c߾}���[n���p�ټ����`�L`�.����0���짺���0t���O,.+��o:��5�Y�z�KW��x�+�wy|��K5� �`� �(�
�tE�1d0�V*������#��i�9c)9N����H��9FB�7�\�@Q��YF4�h��_�`� ���K(��&M�)9�E$W,�i^�l'f��8��6!�b���y7���n�����^�
Ƃ�����ݴM��ĺ��t�J������53i�$Y���p]�~�M�÷�6]/��u��4��0c�`
m`����݂��A0�Y״*�CX@�L0"���^+_)���SΠG�$�"P��W?��\�((�eI�}	��
���%VM�����{+,�����uƚ��R_�j���&6�'�m���/y��F���l[c6W���cf4Cp;�9�}J�!��+t VK1Ʒ�*
;(a�@N	���}L�Ir�_x"!{��LԍF����"TI�����6�R�7�>^^,����J�V\.�g-�����s�T��]�b83D��+�.b�l[[��(��o��#�}t����������7����W�I)�wC�l�Jl��>��'?��DΆ+��_��.�A!�}�bŪ��ܜ),e��5�8�Ź��!�r{�������Ե���G����Om޼6��K����~C���]���=��	,��'�M?�����%�l�5���lc�RG{��M�w��s�����-WL��d��f��ԴhɃ�k*V�*���b���dL�)yM�����<��c:5E��)����l �j4A4N����);���:G����e{�˥J�
t���9z��������w�3�o��N�O�o�MU����	mre���D������'@���?�}�aݚT��k�q���u�]��V��}}�V������i6��D$�J^��V3_������7|��l�&�s=m�;Gv?��D�Zز ��N	�-�_OV�B��[V�Ŋ�4��V�Z�X}����|r��s�K�N�ny�̅[-�� �qv��v�vBhK��P2B~�N%z����;�������O?�xy!��F�Z��Y�{\���'�m]h.KA��4)R��X�`U=aa�/0
�2F�*��|�&x��L����6LO2�l�={�T9iT�����K�.�
�rʗ}x������*��7t̎N�1�1͂��(�޼��_��M�i~�xx���6��}/
�a�n$>H
�:�"9�c�AHL�Vi���?{C��(&�(�S���"�$���m���Y�M�ډC 82dLtE���5�j��=�l�D}�x��Ք� L���`b�1�ɫ,��J��+�[��T�F�ۥ-�b��֭[�b��5�����k_z�0&\ >7�p��"�iӬ��o�F�j>���	t ��C����#��G�ǋ�t<c���'0�w2������YgP�?�&����? +�r ��- ����Q�`/����Ev=s�V���;�G�**'"c�fO �?���U7� ����������<x� ���H���#�|��KM�_$�n�n�3O��n�NS�Mq��S�
8kp���Ơ�|+�r`00 8���	�jӥ��pn�J�[f�Ȼ��A�\\k٥ت�4;\R�3̿����;r�G>M���s��y�����1��Orʖ6���%�jۙ޽{w}n�)L#\�*ev��\,�tہ,�2�.�_�}n���`�WkH����o�k2�MM�����l�M��b�@|�x�t�Ʀ��p���^  ΅�� �w&�2͌Հ\w��I�;a�
� �6����.˥�������=�O�f)���ɞIJoC����bq��a�Hl��!���Pu����_�5�t��-��u��@ݬf�~Bb7�/���Z��Kp
4m�yz�-�ޠ��H��&qV+3Z���XJ7��.�@�/�~��Im5��/FA?�a�#{|3�fR0V$�#)��w#_P�ωs!�C��M/�U,5A��W���ސ̦��8�	�g-7M_�$-�����3uxj����]�ע�Dj�FI{p7�r#�+qS4��r0YZ�n8	��Z�l4եU ����d�1��7_9��x�rooo2�b�*����vw����O�>"������G]��ؖ/�77���#�=�o�??�A�M�P!9{�r���ڲX�-��Xi���>�_�=xMy�0H8Hp�9��~hÆ\��0�
z��K�$��t|V
����Pp���uK��W�ؘM
�Z\��Z
�Z�9;;
4���lo_�^��}�/��/r�T{>���|$;��Дc&///����,-=��}��r�����2����	�X0����L�̈́f�XJ {O44G즁�Y�"�FB7�Ic���B[�Y���1�T�,W,x�7�:о��Qy	�eS�a��P���T
�j�5^�&`�7��b�>|Ty�A�r�?y�=lXӢ���{`bC�i�(;4��=$`B���ߪ1�"�r�'��1�Q��FF+��<�d��崭W�0OW�:���U2�٬���9|I9>�����x��,�dCW�7��t�8��K������V1)Ulp���@�p��\��}�)a��{��l2�^?�w�k�g�<�QK��f�Մ��*��;963��\l�4Q��"�D�Q��ځ�S�@dg{z�T����cO?K��
�)�������|MNw��n:�����oՖ�`NYR�����k�����##�HAd�h$R��r=t�ʯ%��-������*��x%4�}W�3Y�v�� �J��?=;]ZY�U�@Ӻc՝�=�ګ!NB킯�ܗ�Ь.�e�8���@��w�Ug;�Q2@�cv1�Q��0f+�@��Ǌ�H��Nج�EFK;]�/Ey�R���/;'��[�E� q�?�@4�H�4�z�EA�1d���N��	��h���ͱ�yI�VOa5i�ǔb�����B,�w�v��&���cq��c3���#J��H�ˣ�@Z�ݻ��-ѝ������g�����$������s�=⦧�������ٳ�����/.0<G�����?��s�fp����?����E��0rL�^Y�~[*Y<�A�'�2X`�AO�9s"<�A��V�c�S&��= �$�~HK�@����;N�:�l޼y��mП|�ɻ���n@U�ʯ��
��x .��o�_��( O`O�H�������_|�K(a�r�tF� #V�%���eqy����'>�+�(�Oc��L&�Iͩ�M ?߂�C�.��9���p?H�*��V�l�@��PFJ����I�b�s�A�-�a]X��.��A��0b��K�HEL�^��k�r��EdoUp�2_�/^��ב���Hx5��RR1}��&��`0]0��4�����
a��0?�YGߠ�j^�]��?9�!�h���G�!���Y@����O0���Hݶ� �y�w�6lr0�lH�-����Nve'��@b��s��L*�b9AX�f��va�v,�aEP���v��ëij6I�����(a�zE��W$��J�`�'2�1��#����$r�3&J5�W�'�:j*��X�J���*)eF�3˽��T�$��7O�`��!��7aKV�-�ΖY��߭�9�&3\��y�0�'��CO����T	�G���&�,��A,p�'f�3���*�������>yq��T$�Bj�tg�n�v�P`��n}�`���!�r�_j�@W�g�X����������WX�g�ݕcN'��dO����nݸ��R��Ï���\z��cΏ�zk�.�<�+�џ����c/����n�sxxx��G����!�g�6���KY���&�V묶���cE���A�Xވ+�)k���0T.��uyd	����l*��E��:k֠�D0����A�.���=�@���:>w2��%�[PdM�T�3��Y��P.�o��XX�3�	�j�����o<�M��^zl�6mZ�v=��7�Y�}����ˉ������G��Y����c��_��L�����V��{��'kF3�d�dK�d��������26ذ<ޒlX��^`w��1�p��,[�,KVN3ir����]����;�TݮY�}���UW����p���7�-z��Vc��ra��=n�����ƹP"�|&?6�����R&���ъn%2�d�4���:��jw��>�4uD���g��X��c���5��f*LN!��8�i��6��.%���[L���P��J����Z"e���0��av�o�I��I3K�� �����V��B�;�ɏ�_6y�^Q�ND�m��KG1���0�r��e;T�l��ȥ�Sd4��ɐz�;�Q	�Q� �|�]R/���eu��d�J��))n�]	�5��0ʄ뤇'�<K_7al6�c��e;�b�d&��̴�QT݋ȣ����I�Ѡa6c�z��j6��Q��M�۪���c�w�r�[����.���ʝ:q|e~u��]�&�_"����JlǺB����rP�8'<8�n����+��{�}&��ò��n	�N�"�9��h�4��B��� ��H��V��%UKk[ۇ1��~e�؆�\�������v	is����>�Gl��W��="C������+���?^�_�|��:F(.�@��͹����"o"��Ԙ�L�0�&<�c�h;��=R��B�����ȉk��R�t,�e(]���ѕ�ީ���и�/�����#�J\�c���0�a�T�E������v/P?�%*D8��ׄH��޷Ru_��w������8?;G}��\���[oݹs痿�e�	�'�4�d0��k���ǋ���ѭ��H�-���ŋ���!�b���`���/\���s ��x�!�7l�@�w��0�ׁz�0?'�Q1��m)S-.�xlB}��|��k����>������?F����j�X�����b����e� ���_|qjj�̙3
�CO�>O�i���ί�ر�9�,vA�5�'H�� -����~��_���ILxڶH4k����I�n�V[(.X�K��3(l��9e�6�:�n �-M��#�W�D���qF�k�*�o*����q�\�w!\�+�Y!���13$��2ȕY]\,��G���
f8� �e�D.��
����b���PDA`C1c�H��i�!�n>_�w�.yI��&�u�(���-�,���x3U_�^�#�7��3�C��T:�C,7B�;��u��ݟd*��C�oTUx���5I���l]*��A:���ZYY�4q��F��F|$M���>Mm�J��[�D���
�#˰f�O8Hl�MpO�~���Z6m"(M$�`�̚����˘D�z$��Ocq��H$*�U)µ/�tRh6�&����c��/.�7����/��E\��/�e�	��t{�������5��-���e�T����M�v�� �%��(UT}6�񬱿�ǿR*��j7[K��H��Ƿ�M����R�al�veu�ug�t&P�5��R�� �X^3����z��7����o?�k��2�֟;�W �`Q�H���5-[��b	=�]���cZ�Iq55>9R�-.��!�v_u���l�����/�n�妇�����^�"k|lc�e7Z����߻wo�PN���wGJE��q��TƆ��	%NY�=,���hP�u��"�,#�$y(�9�(f!�A`�U+��26:�"I�b���5�,^�^s_,���3��c��i_<$�����-[~�λ���V����_���>��ONl�'9�v��{����W��^� b�����W�7n�������28�v���75��x� �L�ݪ�5�s �J�p�:����"�[�B����J�Ю+�̜?O���g��>~�w�鉅�j��zQ�]�M�Pa�Y�w4jsO@��k�D=�%��]H�O�t���z_e�^��l$M�t�h�;��<�l�40M��I�w�P+a��� 7�H�l��9�f�N�� N��RKۈ<h]���)O�I�lN�v;���z��Gv���rY- \y�AO%:��z��6k�D�
��j���mɭ$� ���:� ��o{��^��g;�:A�ʴ!ĩ�Z w�B:������(̴�p�b���7��TMK5#G�%�V�c�A!��Ҹk&���˃��]ǏOz��bؒ��N�_�Y3���W��"N��捤����� �hfNi�M�aZ���N��4��h6�.���s&�	��mc�5ځ;�Na���?a(��Q�n�B�S��j��5������p��P%`���,��^�1�ԱtSBE�M�T�6k����W�ؾN�7���V!2�8`��l�f�%\���������A����ŵ:�F<�ʂT��6�`8�3�� ��K�8��d�:��bV���J��M�����x��$���̫��>W<f	�K����M���Kq10k�6���_�rV���YZQ�㲔_-W]uU�:/��{��iם�G��� 7S����������7*�=�y����������
���~�̘�A�Xy���m[!�1���2~��й�V%T^Z~A�;�lyS��^h�����'�$a��4f;�K���W5"�P!M�����F�����?�3?�1���m�F��CW�p�/|����b>�噙���ߪ��x Ҝx=�d�,��&��1$Rӄ,c��	��H&-]�+"�ȣ�+�"e_�&�*<ٽ{B��D����$<��Ůg�]�~�2u�UM	$���*�@<I�Ġ	����&�oΊ37F^>�y�~�2�1ے��$�-+HaUSO|�#3L'HOHQ.U������<Z��),��I��� ���o�6S�Zi����]�qx�Ũ�{H��5�G��;eš�|�]l1ZI�R]��=:]�q�y�n� n4�5�
Ӥs����.eg�?Gz�u�真0�m\�G�ZͲ��@G�6���q�G	��>X��N:}����IVt�!ʸ8>lr�=X��K�$���;A�Sˊ<Cư���0r����\�YiY��"��F#>D�|[y�L3��?�L�Nb����������H���b1���и�Q�w�#p�\������Wp	��qŬBtcԠn9�,L�4�����w�1� ���D8��H��`�	��&Q.��Ʒ��-H.��Zz�Ep��%*Q��c�C�����	����(f@�)+��m>�8ݸiP��i@�*��,C7zļ������'�ћH�2��r��N̮lR��<��,ʥ^TϜfH�]J��&��1���Z�dk$Ȱ��ȷ*p�5?2w�΋:�	��̙o|�[�T�J$k������o����5jV\.�/-���|�|��if�E���$R�z�d7�5u�B9��
��@EE*}�9�#X<��0c������:�*ϱ�$�+@:�o�i�1�r̈́��!@���Z��Jd���M���z�;�~׻Ř%Ay���o��گ]C��[wh��;$_>|b��~�{~2����*z��7��W��Ҙ�$:���	�sR�4;V"Ͱ�Z¶a�-J��\2[�:��d�DԵT6���=��w�Ԇq�Ja�o|�g��f.��JKȾ$��c��Zrm!� ��`���H@_�O`�~�oOq��R���2���6VR���vI���#*����pyG��8�E�;Q�BB,�D�:��5T:��iu�AB���⶗S)ؼ�Q�FR2K"���~6t�aN�V��1��t�1�Nk~ ��W+!�$AcSTO��.��RQ*r�E;��juIbt�>DGS	��`b�R���bgex���^�$�0p�г�&Įҁ��=��<=�H�8�M`V+�2R(T��m/�2��u8'>N���c��ka8�B8x�N���;�)Q�黮��ؽ��͞8\��+�����"�#Ǐc��<NQ6iBA��#���#�[,��{o����?k��Mq>�'�{��g��PMo�H�un��r�P#˽�z:��lTW���V����w���+Ϟ=k(�����c�!1/*İD�/V�T��m�^����w��o������K�\m�}��~+��! �R��X��%hu@?��Jp75�Z�����2Z�#���1i��_����*A��J3��VH�g�}+z��Rօx{�8���fRt�g1g\��C��"�c˱��F̽�[�+�l���ҕ�\p��H�J�.�װ�/��z�E����a67L��Ls[	��GG�F�W�����NL���G��_��ԉS��^c�W[�fXK�Rox�l�iӦ����|���W��a�Ȧ^����n��&7ҟ�P� �jK�p��	H�n��r�^S6Q�q�N�)����c�X�����Ŗ��i鹆�`��O�rv�g��\�V_�c_��׾����i�i<t��=��s����U��_#;C.ŧ>�����}[�L�	J!���d:��G"KSg�<9�5;��,M�+��._w������Oe�I�ԝ���c�,�U��f$�ߑ��XM#���Ғ��n��,�u�2�뤃�¤���C|d"F���q�pwpn�ɕ�%�ǈe-D.n�=q�.K�]��L躘%8�ԝ8E'��L��m�͎�z�0嚸֔f̢͐LQ�����i��y�TWƟXt�@|E��1<i �%��E���,�g-m�����Scc���L�����èJ#��q�33�H:ߩ���ڏ؃�_��E�ёQ,����ʝ	B��ؾ}��������ɍd��G���N�N��Pw�����ވIS2
bX�~���w��o��}�GIOm��,-��^��^���a����&V`�a�l��|�رѡq�0��+��I��9���yj��⧥�eV.��X�^6�f�R�����d��q1����lV�^�Rd�Q��q�0$�#.��4�ۢK�C"�\�'G�\@o��+`~��q����s����%�iX횢�ꭎ����Pi.������P�j��.����&ƞ����M��DA����~u}�%��A_c3�}�|�0M8M�z�d�'��h2kc��4�P����J��^}���x��������~����72R6�@(� U�6]uf�n$n��v��o<��'�zfxdL@�/����m۰ ���MS��K8xʥv@��z�1���֢�u��O�V,��Ebc������E�h���f��Iǡ���ܷ(կ�[��' Eo�����vȟ��'7m���o�ϫ�����0������������OLm��9x�4d���ґ3�-� D���󋋵��0.��B�6�a#�P��N��`ۺm7g[�Y�4�g,t�J]�ӆ�R��A�� D@��(�؎���W��K7S��y�B)�iT����`0+�hi��HC����f�� �h���FH���$�Q���d��c����:_1u�h4��Rvjjs*I�P���:��u�'�:�K�qۮ�W��z�VϟZm4�2�.�SP��Cq���j��A)a�m� :�D�4����Rm�kA�5W��}S�4�߬/jZ3JdwOL�:|㬯���,���aRk5�,� �������ͧ��gN�������r�`�Ƥi͟�x��_غN��	�(��H��kwsT�6��4COqؒ���G.����1�ܡ�O0�O;N�
���`ƈ��̶�V�<�u�������J:㇊�H��CQ`(��@��N����2��[�82�,�B*������:v�S�Ι�{���^�~��l)iL�\�x1�
�
	 ������<xem�b=��)�+;7�c�^���ihZv�Db��ňB�^} �ںa�`�*s'Ot�(��̍�������
�:����ލ��'��(�@�?�8��Ls�� �^�h/�5�����^5��jI^C_��U������(���� Ӈ���(]A'\A�uCF=6:�
�fq�@��A*��S+�8���"g�U�����Ɲ#+�~Jj���J<�~=�j��� � �C�0N��r0%0簸q���7�y��R'eC�Qm�3��η@%(j�����?�<�哟�$�"Y���o�3�^�~��5�z�Q/�B�����\\"�ޮ3��<���B�Aj@d���]�B�J�w6?Y�^N%�&S���O�4l����/���3ӿ�˿|~�.U���ٳ�b���{�}�߾!�2؇��!x?�?�5m����\�lQ�qi$�X����,�:/S�\{i[��Z��^�W�8$��iK�:��+^c��E��V|2��(Q�����%+;͑O�٬M�J��I�1�U�]��S!�$JH�DSY�G��A�+�	v�Br�pd�8��y�
��*���֦����/�u�e�v�}zյ7<����8D����Ri��F��#�5�QeRLJ�3'��`>������������NXXX�/6*dkk�[[M��	�H�h#�V�iT���B��m�p����;��\v��������I��wi��W]u�O���O�[�>����ɪ���/;e��{��ez�sg��^����!]F�J�8��fA��� NT�+��m�݆1�|>[Ls�^y��1�W��ݵ{�����S�7��c�F�#,!�8n"����d��� Cq:~y` 3<�Fy�+���P�+F���c!�x��,��M� �����K�hҖ`=g�:x���6УD��88����B�0ו䎴#B�m�E:W
�"n�^Ui��L$G�y�kx`�f,�1��N��Х�<���٪�X�R)�q�ZOZv&Ō|Pe"|�$�ӈ�V��A)�(�^����u�>o�����ڢ�_��{N��Z��^
֫R�ʦH$1M,L?��I�ʅL^�p�<�n�/\���vs�Y����ɩ�?���`!N��ٳ��ᡱO}�S�b�<T*G[��|�U��F����5�	�<����u�m� <�g����[4�Q�.a
�ة�)z�U�]$눃���=#Y��:����u|g(�����É��� ���O��09��◗���ܵ}ˎ+��L�g�Nl�|ۛ�~��J�S��̹T��zm�Xz6[�61l��O����N@@�԰�00�D�o��R#�N�q������ǯ�9������6����I7P�H]�?Ŵ%�9j:�F�Q�� e �T�|IBǧp��$����
+*���2�W�����d��j�)ߩ�t��l�<yzx�ّ6���$-?���|���J{�dRs�j9aM�[K�g��TΥ�sϝ�|1�׏xVѩ��^[(�V���ڨ��4�ō7\���� p��������\�6���jP�m'#_U������	�?r�@k�Ц�Q�2o��{ 1�iU�����,�?�
��o�`o߸+~�o���+�W�[��L�r�[Q`���mh� K(�FF!�V���r�I��u/�X}5����_����-��J(�إ����ѡ��������׎�8jes�����Z*����\�6�9�fmnv���m{w����Q{¿����@�b���{�,Y���r)��}�_����]��w�[�cB-�]ϨQ��-�*�D��z�Z(�!�b5&&����GNb�W	�Iۂiv�L�L,�? �ӯ	b���EU.���	�GUa^CcB�z���ry6&�:M�ۂ#�%���"�u� �1i.�y�H�u�)��ZQ7�	��l���ل��[���	�!x�� R7sؽA�^��J�,�Z��&ej_	no�T�/��:���}�X}��}J"��#��ۤ��J!6��+�����ә��i�
��_�^�;v� Ya�a[���%>��5�=�8?11��~&ǡ��\(��n�E������b�W*M�d�	z<���ň���+p20H��W|���+�8(�����V��%À��G?�;��խ��
��S?�S�L�0�<�W��%��[�^��#��R���?�Ӂ�QJy�I�Zy�m0Y����x�T0��w�*���QQ��)q_�c��E��`�����X�)<�D�����M���\�F˜�c!���op��c.�[642��n��V)��X�_����]���r�r��Z�����©x�M�,(y��:e�}�un�fz�!ӥ��@�R���e�%o�ΝcTѽk����H�>��㸋r�,͹0,�ѣG���7p��nc�,^�u0�X�#G����g�լRx'�%Ԑ�IH��J���(�ԨX����^xa�4����R�!���d��j�BB������o3y[�7�F���9��pI�T�p��?�"�%R���L�t���qT��� ��p�W�6�?���Y���.bJ1�8�8Ų.����H7)�|��]hY�v��E�G��q�C���|r��
�
y������n!�J��D�1k��L��� eɼQ��Z�;'d{�.���sR	��.�3��p��BO"�v��};v���R��C����Y�ō\$ �B14�mC�?M��k:��R�	}7��'t����M�	�X�h5��M~E]�4�kp�\�X7���$�RP�D��HR�)��,�d��ik���
�3gf�N�d�8��R�0>��YY[ܺ}�f⁧�z�ZigrR|{��7���*�7�x�+�~��Ƶb�7���_�z��J��A�<	�Sa@��)='Fa�)��� �v�/`D�W�V?0��a�1�K=~��s7�tY4��%ڳg��>�;�����:����v�P,�Uj��oR(�4�ݸq�����&51�/<rRs�m7|8TU��&2�۪f)��҆ͅ뵣�Q��@i�d�}�kv>�$�F��������v[u=*�a�22	h���n�T��Z�j�HL�}��.��A�Bܴ<R̍Vh�*8�A��A&rEY)�P8�/�0	�
$T�ļ�.��#�U�֖����B�/�`��A��Mmdd�X��Uo$�\*]���k�� ��@,
��~��L)�����Wn�j��@imy%�8�a:a�?����7���b�2�w:�}���ϝ���=q��g�a��hne������(���"�LY=�>-�g*ɉrB��R�x�٥���Ӈ��=k��G�[.w�9��A1g��M��rv����?�H6�;K��?�(�>]�<���abs�'h.-%I!%!������9����-���D�5<2�p�RH�B>?R*=����\�}��N[
YDTS�{D�Lrf''��vr���� ��l��ء�͕�QtCnc�X�N��n�
82���;+>1�e(*�(��H&-�?Q������P��Ԁ����u���I���O�E:@�p���]p�!�&˶��c�B8bA�[.$8v���",�i�h6*��)J�?��S�Q��������q�/l\�b��	&�X�k�]�J6)q?�)��ǬP��5��NV���#�_m�ǩ3���q$$������}%�K벫�;�:_�:�:��F���d����ب!!
F���zd�T��`8x�����(�Τɒ]Z���9��!��R��g��O�N;�}��+}N��+��"a�}/�EЋ>��^��b�9��C�1~�5K�:�QC�]PJw��#dN��~���\sÖ-[���/�s���'"�ZUp>��Ͻ�ݷo�x��&՝B�9�9"UB��(��&v��#S,w�Z2_�re�:���r
����o5ZgP������/�WA�'�[gN��m�b�뇋�]�y�j�Q�&���\�́#ԞT/�����Z��|�^� ��`��3���v�e�婯`·�]�� q%Ά��8sMB^@�aH;wn��S�*����TԊ������-�Rj��C�Rg�`����k�a91JYk3E$H��z��5w�+ 	K���هp�?!J�n")�$�{�F�4<�o��ַ��*×(`��W *��"L�fe	"U�6�ܬ�<��^�j����u��¥0E�:�~�X$�hm��ӄ��:�o��A���B?>0|�mnnn�5[w��T|;���@N�mٖ�S��D����ִ�}���W;���d_0j:��P��?q�ĉ+�o�4�L�f��J���̉%>�V���c۶m�����nmZ�NG�{���N� �`�u3�\��+��MSoխ&E	�%=ߪM��ԓ��j�:�e#�j������`\��V�J��	�ˆ�� 9":X�P��f@�:j`l�:�_緹qAJ�I�zj�ʯ�ʯԴ��+u�HR���ڞ
1��MKS�o����UM3Q�.�Tȩ�f3�4�&���y�wxt��N�a$R&����d��qE�0��� ~xiT�_���3�����ΔMfzf��o���va�$���̦��WOOg�A��8�4�-l(O����ϫw�>|�����3�<��)lA�lt��\�Ӫ�``;�t�����.��|�����l��;I�t��a3VO�y�P�)�8�Q:��	����%XG�@�����#+R�ISj;0*)�2��XU�=2�'!G�9�K^v@y�x���O��������j��5��9��?tУ�{Z�5 `X�f��́�Ly��m������M=�z8E5���ښa%2J�1_+�Ka�#�B4�ҴR������kFdg�B"4sV���i" +���6ku8�#m���<�L�,�M&[�J$U+�d�p@##p�g w�C�5Ҷnc����nLMn�r�Lbx�`�`�w�ht���dT��b.sq����� Đ��a�C~�9�t��lXg��g�txx� gP��}.YT�6�@@�m���7��,�rYPB6��9mf1mi~;m��M���n&�Q�bv�~idh�-7U�g_|al`�L:f�|�񇡙<�T�T~lʪ���I����(����n���I*n�Ԣ�m'����K��w�H�4ݚ����W�����;v��5g�ݲLG7�f�P�����i��^e�h�Beܮ�ͪ�����Se��ϳ��e��0.Gх����ƍ����'O�N�ٸ���칝�vcW<���C[6� t,�-��qB;�!2��Bc���%��
����8<�0g�NC	��*.17i.��B�TW�מ�X*����ғ���D9C�;S�ߊ�j����[B�^�N��E*�eg��)L
M74��A&ӣU[  �j���	O���uGh���i�b������Ə���$�|��è��W۶mtx��h*���t	���(!����FJΊ��7�R�&.E������+FU(殸��=�1��6���s�I���RX~H�Q������}4�������A�����ו�N��P٨�������˞ǚ ��_f��%���Ŋz��ry1NqS���w>CM|`����H��=;v������o�V>~�8�;��/��/��ޣT��
��)!�	:����,qh�N�.}�a��\Z��r��Pz�P�E9��E\#��59�{����6�@n܇��ǃ�A�
�����K��K����D����J����HR7�j�8�[��?����g�>r��;�m�&��}����gfCh�a���4�I�c��������vxti�9U ����b�������k�-�� x]# ޟ���c	�څ��;y�9b[T	#���Md�Խ�O�`.�ڽ{7�<,\(3I	�\6KJԤ>ɍjc�6G��Y�`��炼������%���/�eb*.���rv�� �P��t#�Iۼy3fز(O��k��_�����̤m����a�酱��g�>�k���r�&Ir�c{�N��"ho�s�pwcS%1d ���:�ų����������&.빹A�sp�Ke�P(,�p~�BY�V�һ�()g�S���85�/bx�c�qe�<��Ӑ��;��V�%p�Ǔ��`���܁io}���7�YW��Sq8�	�O�@����5�+]���*;AV��N
�xo���*RH<?�P��Z���&$�nQ ��dM��ͩ�-���s���,K���eJc�/θ�M�	L]]�(�'^�]q��ۭ}U��g/b�f̗@����a#�����@�Rށ�N�(rK`-b}:]�l�i�(�2mC��[���8��yōw`o=��A�顐h��|̲��N���)�mu���%� g���tO����5n�GQ��c�k"y^���YNC�/�r��xK���Ug?#�ɈMf�!Q��z¢����z��a�No&s������ٙc'����[:804d��_y��_�ㆇH�'SŁ��r�A� � Y0E��(\����Wr�_�q۵HR>R�'Y��9�?�?9}a���82x���뮻n��M����s��������?����گ���y�E�����>�سs�g��`��E��N��ԜY���\���(���(9u�`+�_*a��7t�FA�������U{�>���t�����,�,��)ķ.4B��,#Q��$���Z�i��JE:X
a�Bn
���COTb�,�|�oa~Ν��N��a�D���+�!b	���&,����W�ꫯ~��F=��f�Az4p;�L�R���~��h�EAn�aq��P`-�����o�����ka�r��L��T�+X�Q�6��:�Џ�9w�O���_�W7<6p��+�pBM~��8�k��[O<����r���{��?��?,�U<U[�שu�ij���G���k��,��a{d��j��|� �n�U3�ȏͯ�զV�2�U�RV.c`q=���m����CVFI۫m������R�������o�f"kXYR*A-�R���F'���&���BQ��*��ҝ�����$"|��U��hK�UJ��Ir��ab#��CG��[���!��"�sK�ӱ��v�+��ЁC'���֪�����m��R�p���z����6??�0��-[��z�h��mD*��C/ru�Ӎ�ǡiWt#(S��Z�?o��V2�+$%�$0�J)�\�F"1{����®��H�NS=�J�#�e�$v,�Z���Ti�$�����}��3�رc�������I���GF(ÞL�*
|r_�4�_�o�@���&R�Ж��"0sK�Nq,mx��``���!�zɜ������qR~"w!��(����j�=)��mͻ�Y�_Q����+�zq�O�a\�-a����z藳�7Q�{<�䧔�ei>=�_!�D�
B����m{�^w�u����ah�r����L0�Gr�?��?��x������}�c��%�B�וd��XF�#^='���^T��]!zT��Mo���
#��8:��w�[+��-oy�{~���Λ����e�A�[/����?���0��"n��o�����d,�L��E �#W.��o�T|n.>)�(�_q�O�aAKGh�6�1�1#��b�T��q��Ĭ&KC(M�q�n�+�C�ԥ�QǁZ��Q�$!��q�B���5��V<| ND?l�n����n2}*��8����1TB�P{����y�=����s?�s��m�G�N�h���i�T�����+�<~�y��W����+_�
��#�<d�~ꩧ�0�-޽�QX����lٲ��b�/���r_��!Ş={`p��k�[�e�.Su��C��}�S7�L�g(1�k���Ҙd�Ui0	/Ƕ��Ռ)���	�i�x��7�K&�NR9t\�������;žM&�����[GtA;LA:���{[�ͩ%x���{^�]��NF�0��4U��ѣ�{�M@&��V*��U�)P8�m��
<��;�s�����4H �� �iS��fnYZn�ʘ||&�R���W5(���3ew���.E5T�J�J��C���.�db%E� g��N,6MM)/	^�`���1�"6���Y���^K3;ZD��W@��b~������gD%�TK]�Դ�N6���C�LR/����U%r��S�-�UL�,hrn,IcZ��E5�.�a��4��w
ݔ�^�8T�R�ZX�*�X�R�T�`~�$�/{�ڕ�� y~	���c�É�[TF c!aӎLؖӁ��V�z"�[o��M��f�_Cid����,V�];!���k�����2�g`x�������S.cvN�_��_KI��-�cG0�ql�����=���H��Q)ۉ?�B�^�ǩ��Q���t�2�n�4��_���;G�7Ԫ-52G�'<?���%�0�n��G�S�O�}�m�;��GN�����6�?i���9��3���JHy��...BI�ɐ��*�M���a�9?3��ɲ�J������(?����g[pΆ��N�Ө�s�b:_����� ��G#O7�	�PS_	&����ÿ���9v����m���6_}~~�P.H��oT�L���=~�7?�������V0έ'�ہG�/��>~*2塡�����,�Q{���FF:��ҋ1��qr�]�h��t��&]��9���X�<�����-7�6�z�嗟y��Ķ���$5D���dth#!��%�Y^\J���c���[gf[�+g/���ט�������ٽ�nܐ�x�Ё��~�؅�3k)%x��s�sD�p����t�HE������R���*��Rڢ��ιԖjm����_<�rN�<yn͇�k�Kp��ƥu��W�gR�m����~�t��Lme�D�N�̅|�vc�������̥��^]�Ry���W4Þزs�R'v);u-���G���`um[���Z�/��s���}�������TL��n/t�h�Q3�ķ{��}w-Ԕ���?Ymw2�t1���%��@�4�/�@�r�O�ތ�l��/����!fȲ9XB��^pV6m�"�DCW-SwC�22}���	ڵ����	������		N�EB�!�x%c�A3P�v�ߒN=ҟ�Ի,�"M�n3�#��e��eG�wG����h���ZT��Ɉ:E���f�>�̫��U*H��^Z ���b[���}Bn��? ��:F} �~5л���z���#�S���m%�g���t(���r��u�%�*U���/��/�g�b*�e���2��|�Ͱ�\�\:�+�˒��6�փL,Ǧ^��.{�y�1�%F��_�8�!]�������?��������ظ�����L�}�{�?}�Kxw�� �;��/~���۸c6�cPjz۶m������֒!�ۈ2�IA��E,��0�}pZhV��q�[����WBVc�0�I�N�����U�4%1..#�ƤfUf:q�H̘-�o�O��O�ѣGq��Qh��]�bZ��4�U؊�B�l�4y����
�E��v"��[��e7߆	ܱc�Y"M���}N�*|L���#�<��yj��1��M\gC��ĉ�I��g*��v��G}ˏ����o��_������O=��,!�6ML��7\}աC��:LI>���O|�B�6<<q,��y�����|�hgخ���͛7o�8EhN�ei���ߺw�:��s�DR���Yq��V�DRu(�a�ľ�Hr�����Ũ�$�Ɋ�g'���F�z]��5�	����t��ݿ��7nlq�F:Cԓ^�F}��x�R�'�2�;�{�����:��8n]�Pp9+�,%��x�����_�Ë/���]"���n"�bN\�LF�(�(�����Y*Q��m������e32�������gjb;���ZةRl%)	��0"1���NKӈW˅g�P5By��+�ꍖ��H$Wt�#�gH��F���� �d����ƿ��~��5.P�$��q���N1��xrŌ�b�
�B.e�g���UiE��� ">T�T2�Ld*�*�i�&�M�#pJ,n��0����Dt�^+����-�p��6�=2/%�cO��ە�:U���� �lZ��5,Ŵ�,���b�L+������ݲ�Сc����K/��?�=�����C#�I�3�3��,�&�I���o��O�#vޕ>��t�UY�B����,!��#�r�r_�OR{����^�"ƶ��J$
�v�;?��?���Byye-�+LO�h�~�7A|_�8?:>�$|Ue����;~rx�5�L�/n*~���d�3)gH�F�Ԫ��j+�K�Z��َC%�).����j�"��bk&�4�/(R�3Ο?��<7w!���	���W �4SK�I����aAÅ�N�m��F2��x�{�&C�-p�(�B��(�����/�ɗ�ҵ�R���L]E�떽��y�~je�T�1��'NP#���o�������s�p��I�4�{���I8�]ްi�S�ck�3�����epG:�u����cf��-ؙ����Nem��"FU�>�kb�,Uzefevan�m>z����(ه�=�����[mu+sb��Ծ��uڧ�+�++=�z35�����K�j�F O�0ht|��2�������(QS���'[��S�AˑJ\l�mY|�S���I��%����s+=0�L2�'ժ�l�rB�1|%_h�Z����2L 5UP;D�%V^�Zu;�r����T�<6 ,�l��:�Q&�N_��F�y�j���ؘ��7T����o���>Ր�v��6RZ:J�����?��?߽�>zv��?v���_{����=����7���l�o�x��'.�"+�ɕ6R3a���T�(Vˉ��(Pl7��d*S����j��6;V~�����ԙ5�J��W6
î���8��9>sj,Sm��CiP/�fS:�����	Q���(��^�aD�K�I�XmR�)jJ�����̘d�C.U�_L]6wky�13I,=�ng���|"I����5�R��JZ��L��+�UZ*IR��pHh�QFc%��-�Ǐ�BҾ�ƀ�^޷2���޾�SG��ܣ����c.S�j'���zv���W����G1Q/|�q�3�H�e��\X�����~�̄o������Ǉ>�!�SR���w�
(���^��W�B��#�~�ԕ_7��+Sz��*�� ���|��ۿ��(Tϝ;w�$���G~dhh�{�{쩧�ھ};,�W��	�2�u�#�<���~bb����6re�&��Ҝ4��q���B�1ɯMd(0h�h4k��u������Q����Q�V�ږU]��Mg��Ygyդ��t ��YX�ZЦ½jE�>+�:7T��v!I@�}l�c'�)܉)�������ӏ?MD7���hf(X��B��s>#`�F'���Ž*���8��/2>a��N{mϞ=Ǐ�s�Ә�/|�۷��2M�)]r{��c<�� bfoJ%�,Rm�W��#@��M��`ʿ����pV:�+��[k�a��'�$���A�.9H�P�P���t�)�
7�e��$����ժ�e%����$��6�1ʂ`�h���Z���sV"����+���-Ql}|r��M�%im)�[u�2A�3$���N������}v���_{�³��͆��_���x����;�^gu��e}�p��ɧ�=ƶ�2!zTW�-������ݻv�[V�XRj-�<'v �!d1D?�3�Ȱ��g��hXQ�`��1�R�±���Ļ�D1� �Jej����A�.�]c���Z��˱��.��m#ҡZ\? � ^U�p����]��Q� ^[S�z��g�	7۝f:�T��\��m�(a�-%�&ȭX�7��8���Iu\n;�B_ܔ��¶��d���~��3$��("�Oh���nVj_�ңE��B������{�Iq�,(�&0'����BȤS���=��V�
j<�5m#�/��b��Z�..�ω0���D1n>3:6ɻD��ax�d��f�6={~f�+�5>,����p�{��ԩS�B��u�>�pr��XX�I4f&��=�D�'T9k-�3��b�1o{������������p���s��z��&&�1��S�w�}7.<;w�v_\<��KϏm=}�/��*�g�i>����C#�s�R�)���a��,�ڐV)+�JwM�[��y�C$u��\lu��fX/��<b��1x@rq��"�Z�ޤ~5��ٺ�ybd%����Z�{B�����u�:��Lk�Ԛ�*����*�d �������V�%��VZd���V��λ��N�Eq����ŅJ��md�N�੘jp9"
�PK�9��'Ε�S������p��nԚU�0r��L�~�M�)�0�֊���	�tiMӹ�T!Xe�*��1�R������l��5%Y^�B%W^��t�Q�Rm���H��J�߷�͚�Y�CX�^=�M~%�d�ѵZ����O�&�s�v2őD�N�۶�Ņ����X�&M�eS	j�:Dg)�9~�xeiq||r�^�NLNa�^:���S��U�/��W�D�!ݯ"�e��k����L$��g$�U߉��V��2_�ֳO�xŞ��T���O��V���ȥ7�;F��Ω;�n�a��OE��TLsh��v��ȓ�WvLfO���� �!\b��Q6��i"��mߘ�j��B#l�il���
�u#�5~b^:�u��+Ol���XOt�k�_�H��j���hzQ04���:�6A(�`���qB�����"�����(f(T�71��N J�I�;��.��������Z�����6��&��P�	rq5"����R��|���D�E���:}�ri��]H����$K����	�I7��(+i8��D
#y�6��Pz����$5����+��6L�q�Fޒ����/>%^�;^|��|�]w��=r�����i���6͘.��j�}�5�A������x��?99����+���������/}�s��*�d�A�8�\ɑ$���0ȱ�Qh��s�a����%S\(OH�Z��.�3��i��磋-)��P���1(]�M�lN</1X���&�"���r�c0����1�� �İP���#��)�.�B���'�.�sK�b������ƍ:�Дx��8���L:#|��c�p갦Qn\Y�O�y]N�]I�G����$*���3E�<Ɂ����S��I��OD��*[�1X���Q��j��hlr���56J��B�X	��mj���X�ih�sC��
�4д���彺���k��8n�Y�!� �~�����$��m���	�Z�Rz��K�G��L�����U�&��������=��'\����3f@64>eҒ$MEU"��$�Ok�E�z�R���%C���Ԁ�+��l!g}�7�[?�\�A)AəT+�pd���,�8����N��T��Y�仪F"�q�F,�(PR���V�hm�����ض�����GN��&JH;���J8]�	]�E�B/t[�atxfu
��ˇ��Zg�+""�VA��K��^�h��Ҿ~���{"�l��������{Q:i0�]\�6!�|�)�ah'i�Ĥ�[U�����p����Z=jP�G���gs�D2���o�]ӃD2?9�[?��`�U�.2���?��?+�Tů����c�`���'���?	1V�ՏX7HT饵�[�|��>����o��i�S���&����������̅X߯>��}?�6�hթ��z'�}j���<�	���"T��-F�Z�D��
чt�S��Ԧ�������[��tǧދ���O�<�D�0n:Z:���,gU��WתM.Q&�f��)h��r��,�P�#O	�����*��b]aj�g�x%��H����n��Q&�dr�7�qyy�q�7o�Cj3���
��t�[0��k.�r�H[�􊚈��b���6>"�Rٽ�LH���}��r啦k��K��X�u���B��ܸ���Y�?����R��zۄ����m���:O,�=��	L[� ���CM��I�ͯpɕ���(t�B>3���C�/IÂO���V*�r)�����-[�F�0���	J5�̈��i^B6�0��"�HubB�qy5�c�����QaZ*�u�	�Pf�$��Mؤ�J����:��'ℒ��&n��Z�fU[�ժ3�-��녚����L%S�Me���M�&�٨�G:I^U�U���.(;����2�r�233#1)�^�~�F?�]�E�ө�JE!zK&,)��C�(h ���E�c?�0��BH#��U��	u�>]�%Ӵqw���-
)4�6ˑ�4QhD����`~����f�g�a���J/�[M�7f/��<.S}�}��5��ӫ\*\X����d��6���܀��,��	$tN��"��U�e��'�?�a�!��c�a�[�������Ph#aK�s�B���p뭷~�ӟ����
�v!G�o*���хF�\^���gL"�c�^~�e���G�r�̭Vۿ�����s��޿��a�b���={�����+Xz�t���X��!�̎G��0EGypP�1�ŎŽ��6/ϕR���=N�(}���ط4�z;���&@�%)3E>(����|�B��AZ������0U���O�����*�d: F�ZN\q)m3&6�`�P�I�e$2r,�Ν�]Q�ֲ���;�6��_y�5�|K�3E�SJ�)	���@�K��)i���t��^j���������}t�j?n$s�	E���$�\���T6��|`�`>t����_\Z��E�X��E�u�磬7D��GM�T�>��{����xcb�kq?�P�rd��U��(r��|j�ɕ�d��Q�,�n��61����ncD"���xmJ���"�Q"K��r�0�Z7j�/�<p���:>q�xB�v*�i�5n; Ą���l@M���V��6��9��ɏ�BQX��.]D������qۈ�ڹs7顶�����DD�[�P#Yt6	NTT7r����Y~�{=����9*���
�ir����k����D���ǳ��x�J���(Q�е���V�D_����}���P�"!Ү:U��YmX�=�+���Z'eX�����p�m�MϜ��>�܋�>�h�Z�":���:�|����q�ᥞ:uJ ���q�e=�(��%�~��J��n�W����Bz��#�\u�U�}�{ϝ;W*��Q�~ꩻ�z����SG����Ә�0�u����ʓ���{4W��ֻ�  �LIDATh4[9%1]��u=�J{����ۺ��E���J�T �2U����t�SW:�3�(^�jd�1�L�CK�9q���=iR�ۇ���A��M#�����t�s0cCī����{4!�p()�C�S:�
���tQ�� ƕ޼=`Ip [���!b5(�%e�08ѯ4[']3���5u��n�l9��脺]k�ƴU�����Jpy��T
+�-ѝ6<%��n��Vw�m;SH�sz��h�C��WW��̦��p��˙\Zov������~Rb�]^`?��.l���9��;�����B�����g
wNˉ��2k
hȦ��8��/hq����[-j�h�\�K\��\���(�w���\y0?8<��f��ԘA�b�F� D*@�o��{�E��@�v܊�c2J�r�"'2�4�^��dp�������U����Bǧ\Eq2�E��J��S>��(�ǐRe�0_�@����B�>}�Ң���� ]@���TvG)\���?��iӦ�W�i��q�'��1)B��Fև��'Fq��IwF�=�5��#+��HdR�L�����&� ]�٬*[@�R��<;;z��;���^��J��2�;�_��H"!z��)�փ�Zߤ�'̺�.e}������K���J����:}�D�e�A��6#\�D@�3.��f�&%qVC��8d�r�)�0�h<߹k,�g�y�(�X���o��&����~v��={`<~�S��q�U�s�����p��By](�v!�&���~�ea�K�'>�	H���޻��������;`;�+_�5V�8��8p���n?x� $�w��]�V��E�T���R*�J䦰���YRh놞DT�-��M��j]P*�;~ߚƢ�k�I�ׂ��z�#�Z��ά��<,���S��Joq5��^��bsA�����VO�ɯtڲ���_�Q�x� ��*�˘%q��M�F \�ʺ땛���e���c��:qY�,�%�41��ĳ�/�<y�ز���=��K\�K��;�wj�ޠ�!�����=�:~K|��ʾ�*Qa��oT�DM+K%�Z�J�m�'��K�蜻�OOO'2��3�:G��f�TD�5���'���G$��uoLYo��Md0��On�k�s��"���d7�B�����r?�s��0}Ӷ`NI���2s�4l�E���i��E�i��I2�ϴ�����X?�(��>K)�!jq�����������&mJK�Ͼ�Z�>ڑ����n�>����p������$�泃,��N^�Bt�S���?���oP�'��v���iS�T�Ź�G�&C�$

��y
��`ޤe��?UTb���j���l7���-��=�ؕ��%V|���J�1��|�-����8�����BL*4��Q5U���j�$��@Mg��׬T�~���=��o�ر�V#@�����ٳg�������(D0���/'\A��:��n�	Œ���>�k	�A@��۷^�ѣG��7l� 5p�����o�����|�3�+��"�����;�����}-W�Tou����O���`��l��w�����E�#�%/���m涨��	�J�}��	p���iɮ�^�]_m=<�u�J/��V�������r�OS�Q7M�T��+�mVZ��s3V�i6=��M��tb)T���c���X�R�h�4i	�Z�F��`�a^�!��T��#�=�%��sѝC���'�0s&���H#i4(�`a���^���~�c�����~<�!	!!B�P�I��gΙ3'�>��w��V��ݧgF�Ɵ����^�V�_���"	�քh���J0Ҥh#�x�l����!-�(��K0,GaO���2���D��ə��S�X ��Ϛ�����h8b���Z0�p+%0D0*�R�W�ETO��C��G�nţ�Ӏ�����%h�����V���g��\5��>[�>�"���ͪD"!0��Y$��\b��ę�l0M6��r�V���D(�)�<��V�SU񐘚��_���ƥn���U�M� tP����.���\��6�}��AW]l̄qP����<���=܉M�>F<$��s\N����á ��1�-�B��U�nP���`��X��8�5F"��=	�dtTà�u8*߀��{��|���來�{{{YơG3
��Q�N��k��<�#-A@��0`'�jjiT�&A�:F�Ƽ��0� )hN˄��"-��eR����M�5�8�j ��W��j�S��R����%�D��Q�U��W?j���U\�>�W����z!<�8&��NV�H�djg��Z*�0�"��!��c�����ǏkG� T0c�~�az�/.^���={�������jժ�o�t�_��_��Y�Z�W�\kBj���BH�ҥw�y筷���o~����*~�K_��iN���?�;� ��-La\�v-�ͷ.X��ةA�N�$x�����s�l�ۉ,���	 m�В@*f-�Ef�������⦴B�LsTH��H
�(��i̊ܮcZ2�퉧G��T��S�8	͏F<0�a&-p�)�1|C�#6�e5�[��U�&ʭ�G�"b2��k֬�sx��)�id["���x|����ܹs�8��D��&%�~]^Mu��Z��z? �����fM�eflvz��P��K�`̝��#�����o��+v���b>�"e�2��2���A@�Ї�RxuQGx�;��K}}XY�!����d"�b E%|��)�1��,�&�͈2z9�vn �~��˯~l������h"K�E<���&]6'̛
��+ސ]	��4 )XBJkb��%�IH|��(EN�&C$a7TW��"JVqrr^�$���	��iEe=�׭߸`�"����?I�	����MA������ﰓ=� �r��OeK�2#�X��;p+��2��E�Xp�::jhBwG3�&���@�	��xx�s�E�a�
�O`QHN�y9v- YG�Ҍ.����q��l*�*Bf2�(�R��uȪ*�1Z� {�N�d(l{v���aa&�C���UXħE�f9L/W��|�@r�`�j@�<''H|��#	�L2Z�P��b,Az?�����_1�IBYH!h�<E�ǐ_F�R���׉��4I�}����dl�Q1+ 喢��f&̅uSO��P28����*Ƙ��j1d��ki տb�3�#��%�t|1�)XɎ~Ig�zH�V�Z��o `23_��_~������B> ߀�&�$��6I�;�n@5h�I��ey4 ܝ�OM/^ܳa��[n�3S9����?�������A[C#�jjd��o�qh�u�a&��ũ�%���q�W��C���)�,�0q�U�_�����:���ˉ�[�kL���gF��Z@�����D�9�؅=�(�ڤ�-_*a?�h����ֵ�d��簫8����93��> #�R5���d�%�b��\&�=���8ldҒ�pFiA[��ӧ4�7���7I��n�AS��2��w���;ӵ�@s��e�d�/��_Ӹ�>v�Bj��̫�돌N�eL��H�`��{4��&��6K���kY|�)QjuC#�4��3�Q�0������M��S�d��a�������Q4��ڣ���}��S�F�������w*�@���Y=O��$�e`	y�v�eQ�����=Ŏ��l��ccҳ��V3W����Y�ю��ǖ:�ː�{C��}׺bXC����|m�e�	E=Hg�\��o� �!��*��^��+�{���a���q��F_�tA(�YT	sEL��0��-�g�H~ٲe/�D"�]���C��j᫭�(�����>|�u�����[��S�ڐ��s�
p%Yd� �@ڲ�L#�
)?s���T��=�������Laa��U�!G�X���ÉH8���f��Mkj��ر#�*e�4�s�}�'��ڼ�f��tm�f.Uȋ�pjP�d�՜�
^��k��Y��T��	b��J�4WW�\�,�e�5���� *q��c���-�I��AF'{�uuu��kz�p��Ѯ^4��ɧ�zJ�5���]X�����+�����ᓟ��?��?OL�b�qn@Si;�Na���œ$)�C�
�4����a�P�L�ݦR��n�-S.|���]�jG�E@�;v���������ON��W�֭[����U�4����R%�ۍ�@ft���#���J
AX6��bʜ�c�~/G��R����>9,!���b�|i
q�B���49@
Y��Q��ۖ�0���6p.�� e����i��gΜ��u�V@��1��X6
)<�ɠ���J�3�� 93cI�~LB�z��y@���܆m���J�C�e0���E�;X�7������Q?��!u��k�g%ͩN���ŢM�=�ȑ��~�y;���
���'-v����d&31�hEN$ڢ��.�����&6�+/~��u�W8ʵ��'`�:Dt���]���V�����0m�`�W+�	�c���+W�\�����(�?��#�s�U����֎dk#���TR�f��ДK�<��<���%,��< �zHR1}C4d�,T5lYĈ����1�T&W���ǔtװt�E��]'yN%�
�5��P��Xz�.Z�������[n�!���[;}��^{��ð�O�}��Z�+ �&��Gҁ	F� (��~�MM%$_;�di��r��a��պ�n^���X�R�Һį�JmV�.�a����W��T:���&��滄;����#��]yjH�	�uD9�/�J@�����Ě+�m���:�N��L&s������t��$��� CCj���H&=��E@�
����y-�<������l����ZȒ��V�ajX���6���z���ǟ���>�9�}��`Ƨ��V,[�~����d|�LCs��1O���뮻n��]�pM>8<JH���o;&���܌�	�ǩq^E���]"�}��:5�Q{Q����s�A���� ��@�dL:b���V%���8��+H���˪*wĎc�ӓS� �!I��n��)�HD�����	̀)�k�bB�L�������	K�~�BC[���$��"ɈȲ�k�J�h`�xQ�o�T@/��x8'E��bG
AQ1�@��D[z�Z�%��B�X(�-���q'�[��k(Т��^��&�֒��I��@f�[[0��4Ҽ�?�q-EGH�c����ӽ ��r5b�~PR�s�B*�"���C�H$V,�ǧ�l�'�µ.�+³����1��{ȃɒ^<N���J��5�gLz��TD�`a#rV_�iASP(���ɍ��q�r ����l��7���*��.�k�7���25�py�l-u��c`��i�ߡ��I�>������ W(@*䜉a�nQ�h+N���R�"�w0��ѐ����s�jɋ��o��'��K/�4�Ē-��6,[�x��}wϞ=M���!V��kƶƲ@B����*b��id����*�8�?���T	�&>�&�a�Dʿ�q�H��8ն���B&|�h��nL��9�(0����j��E4���wޱ�s 	�^A�o����m�a�୉��/��0��mM���M�`�!�Gg����`�  Z�7500���/�^�����ON�X�1s�����?�k��5�M��(���A�o�TF��VHp����;��`=x�SU��X�<�<�y�05W��K�Q<��1-��Y��)���!�zjp�\�D�Tp������E��?É�˰���!]'u��5k��0�{��� 娸p�Bե"������#,���$����]������I۱��a�(�Fc��֎g�c�U$������>�CZ4��P_%�����rR��{�"�uan�q�KmRO �����5���=�a�?i.r8����0�l�$'�JA�Iϻl^}��t$���LH���u�P�d��g�r&�N�&�;v�E[�]9��i���B0J��@��)y�ᇿ���ƫV~T��k���6��MR�8��N.�|�5(HYdel����<#ɂQ,��U�Y��!b�Py	!��Yd��J)����1
)�>�p
#1&�.�;Lpȗ�sxDV��].��A�ò���w�X�Oe�l��qe��sa,��z��އI�dA9�w,SkEl����9�$K~l��� <e�C~7z8&�����CZ.Uj����Q	�]v�S�AJ3G��F���,�C���]r��M_�B�mI�O����;x�E=qŨoV9��[c�\ٌ$��F�3�h(��/��v�f�s�`���b�z6��fc!���C�(|���9r�e��l�2�U�����\N�X� ��6ߤ�{	0 ����[�^��X���z�iit��b6�S3��Դ��w�r�?��?;w������鹵k׶�����ϯ~6j���h7�������"��~����p%�Șf��3BT�H^��uV�1�j E �Z)��t� �o
�q춵+o��fP�0�������x�M�q?��σ񘘙��Q0��Ç�o8	���ٵkתU+A�<��3�������d<��\����۾mâE�,���}����z����?�'�m]�d��-0]�݉t�9x���>ۿl�֭[MdR�>c�Ⱦ��E�S9���ڈ�Y�l���w��-[�)�ьՑ�*)Aב�6밞��F���-�==�]��r���ތ߂�6�O��F%\Y���={��T���*0R������L	��ƹ�c��Qًդ<|	��iډ��p@@��I�IhQ0�=�����Ą �Z2a�~�2�۵_�������E�����"�>K�I����*|Hd4Ɗ4Ǜ�� �a�HҾ0�̘�X�#�8#ˌ��[��^J�`?�-#wN=�M�K�.K��'kٸ�a��`@�П��SH�aR\��G�0")��D�-̝pM���,�c�c������ܹ���c����!��)�
.N.\�pӆ%===��J0M���҄� q�$nV.K�Q-�e+y��f�&���<<�<�bj ���kz�
�_��z�Q�"��\W��������*��2�r�Z���R��{.3sT���XKKK)�_�~����g��?~<ِ��p��w���w���.[��4�9x��7ߠ�(H�b�T\�0C<��#���}�����~
P��H2���O������7ܰ���X�H��>��O=��c���9SSyP�jc��^���kGG�6ɚxn�� <����wuuI��p2��������X��ӟ~�nF�a�L��>� ngF��f�s ��u��_��W��/�����ڸq#��~�
l6H�퉜w� �d��;� �[� ��n�����O��i�&��`>�P��Yܺu=�dx�ց,���l��ʑ�:Xd�4�v��G�a�G`f.��{h�@��:g�%�u�	��`�l���)5���z4:/fX�aݏ��ߖmdff`#547�������{���i�+��4y���!x4  	XtN���+����%5#(:����εb�|���C_qPcS�d��A6h�[��ё��a�����<i�4j����@xƋk
#�_��C��R�B2s�n �T:[`� '���8^�j��
:�"z�nل��|�IVE*�x� ���~����l��Ud7dHkz�Nr�xE��
%ӎ�׃Q�f�b1m�,�q�������#�]���{Y&��v��l0�<K��x���5�	5���}��Ɲ�����|����E%�����*�	�R����SY���X
"�	���qD����]�8r���q�3��'����0��p�öe�dYb �D��l>���5 �&3f8�2:�ݴtq��I��իW'c����F.-]��������>�w�B�u���fgO��s�G�Ae;�(0��Y/s
�����پ���;�������&�ӟ��g2�2��,R]�@MÆ\�fU2�873����t�u|��N�\o�����*���2���eQ����Zf-ԣ�ڎ��f>�Kks�D�C��䑑�*�l�Pxn���K��}��/}�K ������?��u�WO^\P��{�I@��[��wy��?�����%��.�+LC$�i��o���؃���*BWw�����W��c�ݶm�=�ܳj��e��dr��� {����c�֊U+oݺ�9gG5��3��aP�y����L��`�G��=qat��g�t��L!�v�!+%q���gD�d���y�7Y�T�%�j��%0��㐮�E~�!0n���,��BQh�kg�eI;{�@�\fE���xpUڨx�AlY�Ƨ�KsY��H0"p`�Y���\8�x\4��pRV�L-?(e��k����Cm���1|��J��̔A�A���3�2���j�����T��	Ģ�0=]P#� �熦X1 � �""vש����I���y^N�:Ǭ|��]��DoB���6R�Hl�'\��i�We�&��1�ą�9vG@�H"9<���tH4+�v�4||�8��������R����xY� ��O�G���J\��νɑ;��j��>�X����V�\ϭ���)�<çҶ�FoP���_6���dk�P�v��;��H�FK�g�'a�hqcfv 5L����;�.E
���;;;�%�w�y���b��x��������M7��K ��_��?��?�;p���.�D��� ��P�������o���X@�Cu���G}��[nټa=���6`�X�V�g^�����"HO/��V`�`���J����T�mlPg��9���\���*�dN��o��/�{��K�.���Kp�s�?�;}���3g���v�[ �����I<����^�a�ڵ���_Ϧ�|S�H[],mlDɹ�~��_R�k�	�:ڵ�.�wq��ⷿ��n�4� ᰨ���5K�o���ay6�1X��0�@:�3a��F%	`����o�Td�C�t	%��wDē�u�_�z�H�x�\9/W��2�V���l]X�$RW���<1��Oy�4U�	C�`��/�R�h$��0� `��pm�s^U�>�[&�A?�Ӵ+/x���׿~���ۛz���Zj%��4�~�e[L���މ�AzK:�<�S���gttT
�=�b`�ʕ4χU��eU����|������\��/@�)��T^�C(_	�"�GV���M�y-���= "��Y[��%=�3��`�%.]Wn$Y��<D��J��)���f����va���Ջ����ޝ�s�ҭKc��X\%��GG�eE,��ȫ�t}�X}�0���D��Y��T;<������� �uK�qOr�<�!]�eQ��uM{��65q��������Z���v��tPI��!NbMh�O�ē�\D���=m���K��GHڇ2<����ˈ�ü���)�L�eڅB>Z2�P�a2�OD�������/���jlz��CG���6S�4���^����F">S��D(�Ă� bkj��ƲeG�������:}	�&�R#�ө�7�޽���f�!��֑���o��Kj___8��r�@�Q"b4驚�i��Eu6SG�p8�He��/���)�a��x�S
���)��l�2�:X��'��<0y��-Y�W�)�����ڤ�KwWGQ/����B��śb�DH[�f�,p��������شy�3ϼ�i��`x�������������*�?~6�O<���vm+����S��������}|�?��?]����Y�����﹚�;��)�x\uյtCM!��b|~V�^���^T���*����k��`dL��96G�IP̥��D���V�66T��it��d�D;�sixIh��? Iˆ�t���\�Ż5O�����٫�9�柣���_5���������-���a�O�9�L[g/\���L��#e ��)w5��^��u�-�u�{�U�pW�i�]m>�V�S�#�-\1T��C쒣(�����Ho�c�I���0#?�喲��
�k�''��#��'�$�.[Z4�o�
�~x2ӯ�b�UU"�V�[�Q���jJ`�����	 ��R�[�C�
ҲRd�"%JD�=��/��V�
�+5p)�3p� y��]��4x�BcL���f$	�T�M����c�B��rN�����~��
�RnQ�>��*�̪+DLR����窩M�7���T=���y�ǜ���<$�'�"qD�yBК�P�j���A]�'EL�L&u"��`7�
�qXp�\Y��9�+��S�V�tz�\�������]۶m;��-,�2� �O�9�x�<�?�x�8�x?o�w:�*�h�6��1��u��g>C� ����?hmm}��.���#9�¾}� è@�s�=�۰�@:ͼ�ꫴ6�$hu�^�M6������G�'^��!^vh2���"x�lb���1P�����w�����u�u��ܹ~˖���ƿ�g��L&i9���:��� o0���w�� ���k����G��y晑Kg�g�ko�`�ҥ7n�����*����_�����xb.�w��ݻo)�0�zɒ%�����汖=�BݭV�b揄5<:&��D��Q(fz5�hWqļZ�4�U�fa�F
�r�����Z)���GM-����Ui�U�&��>C�DXM�(�Ey���m�m��t���!��Yy��~]���y�8k/֔~���������|0��8p �F���w�'�A,=�����E ����j�'���U��=<��)1��
��g��\��w�\_o1�ԅ^?�'x�|�r8s��T2t�nX[QA��h�)
���c8L�6Ճ0�*پx43GO>�������e��S96��OM����1 �����]�8�6��,�"|r�J��d�#�&'����Ÿ>�"��B>�*b���{ǫ���@��_f���?�^�j[���yW�>�h=!!R���U� �~j=HN:������G" ��@��sJ�M�T���N�-�� �J@u%���\.�ŒH��k�����������pKOw�����񩉜^h%DYJg3.�[�f�ҥgϞe�$��:G.�|��?Q�=^?�3iE(-Go���2ع�S�< Ƙ���s�|��������1kܺ�����hʁ����(�f�<x�L��pC�,a����^��-4�I���a�%τ��%^��38�aM�/�!�����[�;@e�l�=��O<����}㖝7=��Cw�w��Z�)��*��p6��������*��ͫV����I����� G[��o�~�s�=����7oٶy��ӧ��������˖-��λ׭��z���\��Tv
E�a-wb����w��3gΜ:u*_��?t�@b��8��O�M@�0b^���MT�X��:+��)���H��o���+��	+� #�;G�h0ј��y1��y�C�D<ZRBA�?��Hrٯ?̽V$�_��W����Z~���ȁ��Og�L�4&mY4H���V�_�����׼��k�WW{�Y��g�O�x�(h�Fp04�o��7�;rqƷY��0��k#יĞ6 Rxj�0�/2��+.����&�w��j^?�1����L n7�1����B.e��|��yl'��h#��y�MT$��"&E��e	�8�BԀ��V 6f+�H��+�[��w�}��E�)�,�����>��/�|�Tޫ�bD��H��Y������J���.�Z�.��i>C�v�V��v��W{B����Z��rU.3��x��U����Zz}��K�%$��K	��`��~ ���%��A	)1l������i��6�%�|���omm�������l9;::ڜ�h2q p� r����p�
�����'���{��xcc��cK��*��g�~}��ߞ<�K��`�m��?D�{O�zzz�9��=���i���J]'�T��Թ��.�JK]�S�/�*Px��1Z�?�Ƿnݺ{M�cp�,?�FuBN;7����s>A__��w/\���#�����8[o���w�~���~F�~���۶oݺ�|�駟nlj��Z�p�~��]�v���Ǐ�����a�r�� `Ҧ��P($ia�
.�,�[0ԂQ�Z�eHP�g��^�I�Ϫ�A#a�G��q���\�1p��ysm�~����2^}�W�Q�~]C��-�|X ���%��q^��)�'6�)���Ơ��l��a�S9���W�n�+��{����y�	�}���{�!I�ݫ�Lm��]��O�ȱ�5],���0�#XE�h��[�f�?_�K�|Qi��&8��+f�A�e@����OY���8屵�	1�~5�8�*��(�J8� ��iÊ�W2)�&��<BHD$����	��B��v������=��Sz:����a����~PZ�9�s�-!�LDm��9�-�0�!y�e��ABm��faj�:��y��,*�4{��z��M�\�{`��Ѩ��D0<�$Twq�$��� ������;=�	�na�Hlu,���1��!,�`��I��z���x2��Һ^vl���³tǱi�8I	����4���^v���K'����y�իW$7��ڹ������dS��U8�q@W�r���X�a-$v�5 F�?y�Y�6nܸs�&���g���}�����%?L����b�d �-�C��S3�ĥ�3��R9�f�lv:%3�VM�,V渒Y4��&R�鑆:x��p��L����lk��֏ݵ|�fP�w�����H�����������m�:�&���.[�a�Ʈ7��g�vM�k6m�t���KW�?{A�#'N�y��=�/�����#���_��qp���'�O�<sq�������MAذ�`ܞ��Ǧӭ�I�����J8s�)<������i�L��(��Kec.��D�$S +%ނp����Q �`�k�ty�E���<���q��W[L��x���G�C��1s���&p�8'���>g����
���)B���b�N5�|���|���DMMg�<'�����a�����􌳺��R�;?�k���j�k������R��F	���JQ?�ё�LJBH�,UH~�K�T<�������}T;���sǢ������8��O�Q��R<R��Kkk+���+�v���
Fj�P�2@*G��H�-���ҁ^��C�4v�FT�u1y@LC�u�fC�N�ǌ�	��㍀�T%
kF7	"D�D};[ۄߎŜWc�I*��4릂�胜\iWk��f�Wگ��?�U�Ts'�'��ZUe��)O\�A뤫vE����넽� M�ꂉ���r��bM���d<$��H�W�����b���[�_�S�C%�9{�lwK�o
�׆�B�%�h��+o�L��c��.�J��F�*��'�GXz rb.͞;s��3�<s뭷�22k�~��}���_���3�`f��T	��`
soo���$���5��P�1��4I=��!A�K^=BOSC��br'���p�'N</{7�x#�����m�������?w}��yEY��hQ��{�?�����[o}�/>w�� ~�v��_��g����#��¼����<��\�b�M7m�]y���ѣGA,AV��_�ez����ڑ� ���P��t���$wh0RHCG��V��*��_=�,o^=Q�u���Ц%X{����P�]�:��ICU�9^�P]���=�_Wd}���=2�Z���O�@�Ф�~Ս�t+Suz  �4O:/�v}C��_=�`�
��p���?��+�E��*k��ւ�/S#��CP]����lm�ߗEԱCKS+�h'�~�����=��U���s"Q�-�l:�`$�,�'Z�hsq%$�r~��z�[F6Ҝ6�S�6�b�1-��LP�8�=,>Σ����;��L|6�J�U,�M@[��Y����ߵ-�f�1�Vol�Ɣ�L��T��� ��y/v�ă���	I;�w|�uN&���Z�(��ޒ�[������y�j#F���Nw2[ɘ��)����N]�Щm�I�5�E뭨q�U���C�a�*�:{�C�%m��n�eHMXf��T�δE�l��9"�(2 #L����b&W`%-o�`´d�l1۝l�+\��5f@��� (�������3�FD	�Q3{xj.
;6�;0�sYt�|�$g���g�rI/����޴n5�u�M�DK`���ϽyԜ+-I4b�[9���}�-�1CA�����D!�ܜ�J��{��D��9c�
ᦲ\�����I�\������{�]�ۇm3�w�}7@��}��U������` p�03�߿�>�ď�S��X�L��E�����c�I�uK��}�=����cA��򘞞����f.��o~����8r��P.��1������O_�L�8�����d�E�����#rK�Y}Ta�,�!�ts�x��y�ʉj���48�؎k�$��aj��>=�c����+�േP-��)��;���;?����G�j�1�N�ā4�a(��<�T�@aHk�(*�cȵ舘�M���9򫴉TYVJi.���j�W�Q�����o�W�]�ڜ�$0�L�h����Jx��r"�"�����MA&�S�Cr	����*����}l���y��&�Ȳ@[7Ԁ'l�R΢�ڞ��.F�)Q�K�ٕ"s��Bҿ��m�FY��!Z�ҟ[��g(�'��0�'
SSS��D�v��$<�6�V �d0tn�H-zR�� 8�\�g�g���q�_���_cx&ǹ�\���VOt}:U�-�͕!�J�W-�0��!��!9L���ao�L�Cօd�T>Vm�K�e��L;`hWO��	D�H���	Oj8���cւ����|F�}|^M��a�a�E"	���Ľ!3C"^4^�L ˥�A�����;;;�~�m�q��^��G"5hoȝ	�p��,X���\����j��N���L��%��+ Ͳ����{籚!����,�(E�X����ߴ���CX� �~V`ll�36��&&&��0BR���R���>=���H>,��������й1Zր$�$��rU�������yD4���� ��p��ŋ'�h�AP�y$����J��N�Di�)&�RH��G�F�r�NO�����	/0��_��ɏы�u��C����z߫P�-�W��.W���IL�楔�ՆB$�@\�z��f�~�r�m�+�ϓ`@M}׻)z��W��iy�u���D�AA�*
��Z����I�=�����鑿y��@��I��(�D�{��mtON��&W�'I��p���+��ND��A�`޷��۷19e�u|<�r�P%��6S�Ǹ��0����Q�Z���AI��k����lHģ?04�$aH�͚n8�htr6%��<�c\���
�_7�#�.00�}�T.�J�x>���ga-�e�: � &I���	�c-��8@��T����l�@��$"�B!��2u߳�n�R>�V��k��NJ�r!7��L=;+�LCS2�2�ç�c�XP`bKK,�)��Υg1�㤳�Bi��%��\:�ʲ	n��ѐA�A5$$q�4� EBj4K�g�y���LQѴ�Y����f�s�p4�T0��638��ؘf0:\2��d���Di�ꍌ;Z����_=4�s�"W�nA�"�Q�3�'�
�Hr�iڂm�����;ŗJ�g�%0'˧��t>Ov���ww5vu�<���͡�Ԕ�5�9�a/�,�f������S��L6�H0�u�xidl�K���xwPv!�"����p��`�G*����T.�� ��UYּ61��L�5��LP�(j��t�!�]� 00���3�h8j�т�dg�5˰�d	4��۶�i�#m��� �'U�9�k��;fy6����h����e��:�N$¤U�)k��H ����h4�ϸ9�7�Ţ��waՒ�!�udҎ =�����"Q~j� ����`LI'���L�F� ;�� �|1�]V�])�j�X�"1,�d�����X8�S����Sc ���3=d՞���f%,ǋ�i9���lz��8�D<e	�fǱś�z����a	X�-�쵲^�PU ��x-�'O�
׌�"�ic0P,�l��n@�����g�tM�z:0䄺 ��M)�g0�BX�<`�����*�e3�
V���T
F��);1��X:W��D�:�`(B�����L
��s�nEb� ����T�M$d%�J	���E|E�s�R};PuXM)�\I�K�<6�J��xn.�!XG�?��^�Al���Sbd�-j1Ib9���^�)6���4�P2�K��|��A�A��әﱥ�E��1��������E��*{�9�%��$�/W�E�\�$З�Ib�mJ�z������r�q,��%R�[����Յ^h�&et�)s �Qf.�#@Vry����_� �M�D��X���G1R$�[��+�����🪆}h���47�:PF�M�X�]&�>L��)�h�z W�\	�l���a�8}�������%0~0-��N&�;�2V&�<� �#���ݢ�N�$�7������ s@��(p�� �R^�è<L���q��WW�^�_��׿~�M7�?~�0G��1�����T�u�$y�ңʔ=%ѰB�RG�qGׂ��_~9��w�ۘ�-�*SE��H�C���\�R[�j ������899����4�gi2>����,qKc&_\°o�z0���	�� <�9f˖-�;�]��
*a<�	D�
���UX+��_5ϋ����κ��NO#l�����0�Z�Eƙup���bh�H
(��E���m���k	+c2N	F���`��"$oj;�q�����i%���:^E�!� �#;��Q��yй���S6,��H�``�M���I�[��Ԯ��WV���疱�v�QaJ��F`�#�h�T�}�`ʅ�$�$��nq�]&�2�һ��+:�0r����u��>�TJ�v@�AtUI&�I�&F����H��D	ۻ�pP��`Wj����6'���.b��!�Nz�ؓKa��Q�aeyz�Fw1HH,!q�F�3��
MlP���0��"��oS� �r<� �	O�j��V8ц�*a����p�PB__��Y��r�6��Φ�x��f�e��3JE�[-��L�<&���*D�j���bc �o��T?�`�&�s��Ŷ9,���?��	�<�@�9`��*f����[E�$g�pG�,���ѽ w-�l�L�?E2x|��1�g���D	�ur�"��LDI�R��K�,�V���vP�yC�E��I9dX�x"��.`�Y�TLö�E���K4'�Z2R|�d��<���|�a3�<@<�E&DY`�*�XD>.�xq��9���,�1 d'G�B�������l+����Q|o��>��ӧ���[��(:z2C
�ͩ�m�L�)�Z�e%��E��e����< �O)b�wu��9w�Y�̠*���s�p;r߳l.=�B��<'Kb)�RPT���3s�I"�V>cD���0�����\��	vk�#H,�@���a��I+���5�-��� 3n@�Tte�1K`vx1	LIL��bFoP8՗Fi��lP����N66g���I�B��x6�*<�/�r��֤��ښ�6�5Mi�&*Ō�0��2>}!�@����R��ok����É"�TUH%j8�b���`���lJBT�,Q�>����!�G�����`� �-1d̚)���H!�X�h_ɒg*m�^�����m�i�� ʖ��Ŵ\;=;��x��2���h�e$/a��G#e�nH$�4ɴ��L���%18��I ���X ��c���8�H�s�tF�-�a~���!��q>]3Cϯ�j���g-��9q�u��!�=���ǵ�[6n\�r���c�bA-��(1�����;�/���P2��a�fQŃgKbʪ�d����XL�[F.o{�*�~*Δ4�S+�14~2�v�n,��0�PɉB��w�66����\T���榊M O�W.�]xz���#���a�����H�L�Q1��Eۏ�ε�%8gb�����_:χC2�հb�;�`n�n��N6%M�-d���%�S��r�=��_��Ģ�b1x�w�b>�"�p�*O����LX��SN�olWEϦ;��a���&Z:;�n�KN"jX6o��,C����dK�EM�Z,�`m�"��n	  6�� %�]rXUP�POɓ��d>���R�XP~k���n��p(�Bh�W������0�Z��T[6W�#�?�Ab������*�Q���T�ĉ�֪(�^�������?x�(}���v�Z�t%>v�ؑ���u@�X�:\Z��b!m͚5�=] c�����ʪ�� �=����~�Om�bA����g�f<hX�-��Bo�=�w�ihl�a��W�\�ti(�_��*7hoo/"t3[.\���w��{�zdǎ�M��>j�C�Tzppp��� @���{)��d�p�˿x����%?~FX�M7~��Ɔ��'��Hp=���H8v�747��gN�8r����E������,&ΦA���2��T��k��ݻ����?5s	�2ɶ�[^�d�}�~lϞ=��c߆[+�1��6���8S�N�Ĥ_�F3�~�����K|�G?���� �Cc>n^�
���ɓ'O?([&��.6���w,,6�	����$p0K��7o��׷ V��ޣ4���;�֔�3g�<�����P��B��QN R��l3�]��p�?���c�= �	I�ڹsg��婧���+Uа��nH�{>M�;>�F]�:�����G.���el)�Ү]�:�;������^~뽋/��3#hAJ����:���
[O��W(��Z*� �M���=�\��#Ju�K�.�X����}���	$�݃'h��lEk�I��)޸�ƣ��F��m[��x~���a  ������K�1�c`�QEq���@�ʄ��p��Y�_7L�V��N��(�7����+�ʱX��W�������Mx��Z{{;�,��m7�����{@�s%�-���r��6I���a��b�C����0�lj��薵k��l4����=���O>�{���ߩg JT?��?�)�-����ܲ���[�tF��&����o�O�u��^z�塡!�#Xz`��O=�C𤻺:@��R4I:_I;|�,	�Ei�9���/���}�;��Z&z��X4I�a�[]�r5�#X,��hSӓO>9>=~�­����W_}u��Չ>z�"Qh�/�_���~Jө9X�3'���^���^�;�8���|��wϞ<��¾N�[�U<�%=������'Y������GK@Kz�N^��}�Sڄ��	#&��F`icBL��e���{��b�����!0W'�CQ[<�4%C���0��M��{v���iP��oؾ}����E�M�Dރ%/��������,,ލ�o���9<l���O��]����^�'z	c���׬\h����_����=�5b1�ĩ��_�]>m]�h��ESS�_��/~K���;����1�ujj��ջa���t�U���vl���5�2���]nݸ�0S	Y
�����ܔ�8f��T�k�'W,�_�0�����o��"�+w�~{ggg8��vq�UȦ3yN�%�Tu�,q� 3k�:��&B�QMs���n�{�����~��& ���I�Ֆ��P�q*��F�dy�,A�Q(�8시+q��ga��[��#��`��ĉ����j���{W,��m��+6�}�G?==2T�Kg�9���)�0\�]���p�6�7�)�e7�|�-&"�=>x�s��#���O}얠̔r̲�� =��3VDf�Tk9��4��Vflp=S7|7"r���������oX؟���/~��8��`C��pӧ?�p�b^~�i;���3�P��"��%��زH��)~Y��R9[��-�o�yՉ��~=,����x��{�,��dY��x������l:D��-�D�z��7�����`,��9�Q�l�k�؎���X+��O=���@P�v���+�f��͛�>�쳧G��:�ʳ��\��$�*��WJ�LT�>q׶e�]x�>�M�p{3�����\B�^b&&�c�sE=��OYT0WEN,qn|8�/�l9��)6�T��v��v�dG�Eab�fPdz�nޜ:�[��/���Ǚ#�m�� ��Lvo]ӗ0fA��!-�6䘲�32�`��Ͽ���hP�p%�=�k�@{�O<�s]�J6���-'9�dbl��3�L��}�[�y�e1��4�ln�iU��������olm�~���2�LL�ݰ���[:��!,�
}��,����K��^��~���ʠI2�<�_�&l۔92�S���a7,����n�0%��~��E�̠����]��0��l��O_4rs���l^i�3o�y�P�	$��,�\�w����՞eѦL���ɾ�L�!��^��մ< ��v�eƎ��k|�AE�J��U����\��˳��O�kt4���@R$E��ÓDI�2��xwٯR�)P�<42�w���)�M�[�n�l*����r�w�4%�G`G����L����~4���O|,�ѣG����lH�!Rz� �m�z�d��w ׬Y� >9;��z�]w�*yp)�w�,ri�����/�~���C�ɾ��x�����P�o�a��E ޭ�q w�;�����-��⋠�7mXm��PpYU��D� ϝ;wahL�ljꡇ*X�W^��0�F6$5�c^�]���ŋa�fg��69r�h��ݛ7/}��wN;�w`�p�s?�9FU�`�s:�%��^x��������a��a�W�X����R��ն߽n�ҥ4�����		�O)�iQ}K��J�O�%	�.��1Ɯ�/�VK����7��w�������u�`���b��H�%,^pH��ټ,i׃�h`A������D>�,]���0��|��J��?��G�o� �R����ڠlCSA��|f�j$����C��e�3�,x0Kp�{�T�]�8�K	~���>lS`>�Fp�`�A����W^�/�^������^O� p��,��R����~���:�	3O;�8�	S
�G���[~v��c�=vÎ�?���uM�����zu��?����/����a�C�<(������wܸe����Ny������x!�^-[�l��4�
gϞ�ؼ`a7(�P�3�f�D(qV	$���nܻ�������W�,]S�����X
6��C�o�������ڵ��჏>�h������ژ�1�~������/L;L�����t��杻nܱ68Ӱ@��_���GFF/[}�]w�ڹ��w�>��σ�r����in���?��O�:U��5?l׮���<���G�{����;~x�������-l�#����	^z�%<�S�l���. �«�<	&m���w�\r����ڽ�� u0��u��?�M��JI�}����J�^��0�m�6�ʁ* a��&�4p"=;�sJr` z����o��2I_W����F��^�++!t2E�����?�����u�G`��8t>�ۋ���ȥ�z@� TV��f�*�����뻢+b�7�uXi�<��E�s��3�|aIP�}�Y=K?�DY7�'X�Xطp���{�A%�H�Jh@������+�^�%��UΗ
�\fƒ�|=}�uS��{� �=zhoGkr�������Λ��R0���=��,�OD$E��,p�t;� X�������İ��>-l��e&3=�&�mu��a����xPs�Y��ʍ�/��/���;��lgLs�)�s�����;�Y�B`v�B:��ن�ptv������[��	*� 
en
�\c%�,t��%'ƧF��hHl��g���5h"36tꭗ��������ɘ�Z��j��herH(J���D�,*�DW��J�����XXr<����7�8| Mv���ͺ��W�_O63|�3IV�Gԇ��'�)�$�t�`�M+�lX�3>�jD�����(_)>{z���_���K �G��;2��MPϤs���c4�**`��`�px��Vɛ9
�5��O0eͽ��s���/?�N�E�3=ٱ�����C��i���� ,9��-fF/ߺuˢ�NUdFΟi�h^�����^	Śc���L^�B��xL��d8��Z4Jl��t�9�i���\����+t�Ϟikk�{����Rjr4�m�kV,�ۇ�.�障Ńh ���i�s٬�*L0i��͈�H�u�Bf��˫�.�ۻ����0��3�3����1ۣ��P��������ݹ�A)#J_&y�
[�]Ry$HD���̊���75u	�b-!��������?���3����<9�������z��y�*`H$[,�p�Vɷ��`Ex3�31� �9ו�D��esӚ$92�����c���ѓkzz::#Jw,�첗a���O��a[�
i��Q�KLqb���}'΍��M&� l�f*��� "����|���|z��;G/\Lÿ��z���������A��h����6�E��~����q�r~���D�"��Iލx������M��=](I�kV8�a̩���?t��|�֬^Գ�{"��L�t<K̦��]���Й����֧����|̿]f4EeL+�i���߼���;��������DoNu+Wu΍ЍF�` �L��%��$Kֳ=�l/{<��[O����z^�=��%[�G%Q)Q�E$H�4�t���Օ����sA�f�y?�K��V����s����������BD�\�f�ń�,Sd=�H�/��l���+��Uh�o?p���֎�&Ϫ�B�>v�r��<���j�bS�oq���qʫ�}M��:&�����~I�|�p���Sӗ�;/t���a7�i�Y!�0ba�9p�hKb�3&�[����{gg'bX2Jџ����}�[ߒ� ����ދ��ÇGqrz�<ֶ��z8�k��
F�y��r���Y{��Ϝ",��p;8O,������=�F��{���.�?�dqv�'�a#�Yz����;�#����;Z[q����߅[F�u���E���ۿ��xԏ~��>�x.�������O�n�1��g�gDUI�9���� �T������^�	@���z#߲k��T.��@`ak�w�y��7�a���.���g��I�9$�4$B�y���bJ�E`@�^xA����e�rˁma`G�eG�a:���.�ffK��3�D�ֆ����{7��8���Sx�����$�w�~����i���%N�c��+!>�&?�T�&B+h/v���E��b�Gr�?��?�XD��C�̒D)�ީ:!����U!l"�������ۣ?������[>qZ7=�F��0�������Im�����,�������jۦ������J���#�ܹPmĨ��cMM�+
y��_����Dx������Z5Z;M�"�N�����9s�ؙs0�7�6<�hjHC��6�W�%����A]�Y��'h��gsK
��tFW)��ĳ��'?��������E��1������~���R��}���K�N��G"w�yg{R���B	�������^8��gQ�XS4�裏6f��|��o����?����)�n�>v.hL�=��~�*Ɖ�/.�2��Ojd+���R)����Ak`�o���?���;p�@��\_��W֢��z</���К���re�T�������ѣG�6�Ȗw�ĉ��ka�<fӋu��Mce#-�4��X
kM�BPy���m��/���AO��?{���w �}v��-�����t�䅑��C���^x���MRk��-�l�x����N���uE���橢�I&�بn۶�!E]L�l��fg����|�_$F[�úLL�c��װ<����M$®�z�놿�/��Mu}��4?�GXW(EQM�D͆�j]W����Z���Ou'd�`�NJx�$'���9�am^TVbCi��U�n�����eA���@�;�l�'i�e�q���@8��-����[�3�k�z�,�~2�R&��+�iʤ$Mݱu����k����bp��ƷS���tuBEvx�9Ӑ_\�q�
��am/f6�M��m��F�4����_�p��_I���X��vo��&���=����.]�UÀOR�x��5������-$��J��mm�������jɌ&\>ުU2+�+����"��a�[�l~�����<62B͍gn.��!�T:�s�,F`'**�i<Sjף��ܺ,	A���נ�#K�l<�֍>�s�{�;�
Q:8S�p^`F#E�Լ3���3V;`@ߡ"�R��}�ލf��7o��S+m�x�p�{�f�k7A%���S��_z�%)V݈U�����J��&�qC;v�}jr�����G���k޸t�5�>��S�o�±��dԬ,��qe���7�\Hn�����iJ6�F�rym���斕%o]�Z*���vl��������@nqfa~6�Iu��O��y*��*9�7� [�t�F�T���A�!������E��[.�nݷ��7��V�?{�0����?p�w�qס�|�+�&��Y16~B�����jͭ�{�;�Jc.����~C�MC]�ە0�h��T��d����Z]���M�%n���O|�R~�3W2�d�#X�1j_�f^R`����xirx߾}C[7�y]_[cV�����<y�=U�4�6l\���}���鉆�&����)�"jD!�����D:k;��wn�ʵu�����0�����_=wf���$����_:}�*#�Yس}�K--���W��y�u��MEZ����6dI��՚۽���SdY\�W�񝗎�r�P��׿q��ح�����;���߷f��?��?�.���f��j��D]2�պ��5���j�К�j@F��=y����ӹW$b��_��U��{�����v����}j��Y�8]R5Iuj6 >����_�J��L^�gu�j������lX����{�V��^{��RٷYQ���|,�lji-��7���&�=t��^��*�\LD⁇����|P���E���cæ���/s�:���_�&-J�l��p�*��O��q��x$E������2�I�"󿹽�~a�fBX��X��~2=���b��4��9p|VXD;�a���I��3�9�X��L	� �e�� �P�>�j�Z�r�Hlh6f₅R	(�ŗ~�����>�2�x9� E$=>#� � ���g~�fbb��^�x��>���A�q��ׯ���ܹ�T�LOO��?�����A���o|�ckmm��l@�0gHa׮]PZ ��o~��/�+@Shh�D�QӲL,/Qz���4e�W+=�.,�ʋ/.,,���|֫�yd�ZY5f��ك�"���|���<Q��k:�(Ϸ^��?�S��|��0D7��J3�hz�߾��NU#��q �S�.��VV'q� ����[����]*�PU��DB��$�1�S�v<blݺ���p$�i�<{v�`��)�Uk7'>��;zH���]K����ysi�����˰�˶< ��������������h,��rEǬ66P��+2�π��r��m�2 I��r��?�c�X���=w7biV,������S��b��7E9�5��T�D��f���vw74�s��1��p��G?��?�A��ׁtax���D=`�XW�8��T�
�D�}�@\�DX�G=4:��ўxⳟ��cG�7׫!N��Ttoi����_#w������Y%M���͍��+�N�?���x�� P�g�yFis��XC!QҨޘ-
�	�t�b�P��_N��}��_�={V��_��+�
b�l��q�މ)���')!;�����+��J	���4�b$�;�9��AI6�����%�������"��L���'O���s����m�]��r{�q�N�	2`��Ә�Px��	���N�>�����]1����!�ձv�?������m����W�@S�BU ���xv\Dӈ����#�M�ъ��K�Ƈ�6"��1S�n�|�\�C\�aͪ9rd.7�{��{���蕫���V��a
���]�65E{���/����cB����o��%+�.γ�a�&��Q��)X�:/���+�܀�;�%����Ԡ�!�<'GF��H$�%��D�P��Cɪ�5�Y�F)"���Ay(�W�4+�B�L"����ڵ����W�5�bQ��j����uˉD���?�⥗^R��^q����}6	���V��<�gM���p��ҋTb�H�f,�� T�|�j�^���6w5_\Y^5��iii��z�嗇v�M&���AĶ�ׯ�T��efj�[L|�ۆ�SS�5�㽓g�7nٰy�w�S�9X3A3�,����%r]
��Rͩ9�j����˯Ur$	Ϙhl.�����1�(������%��w�?�e���׿����uk�%3�?R���5��^y�rX[&A*[���-*�nF>�ZU����!#XI�鞎�+�.RR�Jm�әl�)�n��W��:?>V����5g1�蛹"�_�I��GhC�.d������K��G�@ܖe:�i�og�Mzxۖ�_��w�lR*UaO��,}f�,�.�9:=�v?Hp�=��V,���-/��j�u�m=}-�w�}wW"	����'O<��� z�0s}�y�F�TD���{vt$�MV<��7xG��w�������pcvb�ݸy`���J��_%� ��|�rz�%N�ΞH�z6���ƔU.�\,Kh&�]�����7n��s^��/����n�]�}���2�~e�R�dLRJzĨ�RE�W��s)R�f�T�"�ڵ��+e�:_��uv��ݻ��Zi��m[�w9���s�О@11ω8'��H�ju*&�y"u��W�i���J��wwt�S�s�-L^�������}�~׏�y���+�ʘq���k��|�Lۉ��vr:is�X�r�t��I3�����3�P|��c6����}�6��o���?L�әd6_�V��r��މ�w�5�nJ7$N��v����m�d�Z�b>���y~n�,FO�\������>�����s�:׮�G{�o���~����~���?��?ھ�;��iTS��<�:_+��ܘ�%��,˾xbxS�Ə��ѩ+S'�8��w�[�f���5��{-A_�q�%����O>��C�<^�U.��W���í��O^��b �k7lnl~����0�*�^�r��ko��in�r8.w��ɩ��s9݈	F�aa�I%g�*�ji��T����^��|=1�#Z��M�κaJ�
U�|u��Ç�bD��ɂ�ϖ����2q��>|�\����j�J���\��3�������핕b}@F���4t�&�q�a�<'y0�R�aP[�ŶnJ�(U��������B� s��.�1��hy��|�J1�Y$��w�����m�X� � C	�G��%��ji&��vmSç?M%��ѣ'�z뭹�9��fv�uaT�F'�u7�l=��a ���xF �o}�[W.]���㎏��Tf̘s0�{�����
���:#i�s���1-���g�<�60/.H���D����Oʪ�㝾M}MM�/ޣ���N�ku������-lY�jKS��ap�3�~q����Ǣ�zX��{�ǜ������痿����@7���llhhhfq婧���!L���ry}��ۘ%.���#��{38884407Wz�w&&&���+�Χ?��e��}L�Wd���J�ĉ#c󘥰8����(��1#�%�����o#�x��C����[��m���;����
MH�5��%�0 ��2���T�ۼf�޽�e�������oA��n��e��W_���?�@�QL ��6&����q�]��e�S!	��xT�ZN�Azz���cq�ba�ӟ�����oj2>�� ����x�ps��jR�Y��=a�<vY<]%����Ϳ�[H5,��K���]�Q��nnHB�s���ťW_}�F���L��릟*?+T���=��ѳ'������'�ή�\k�DL���.-#���l32Q���댧���Tj��,�����i�[Q����7#�Ƴ���ݝy��u`X<2��[6vv�+
��_�"쒆1C�(Q�����0��Ǐwv��w��������߿�O��O Pj�x1�� o��/����[)R��K�%H�<f~��l���/���6o���ߵ��]�|y����4E�SC$���M'(Խ�޻�J����/BƢ�����E ��v)`-7��q� fszb�z�0-a��%�˘������!��ǿ��o�S9Uˑ!�4̤!�EL��'�;3��˿�Kh�Tn��Z��t��O~��#�<�ooo�4bQ\���e�0����/����I�
�!�x�p�G��͚oϳ\�dU�IZT	y��25��-�EII>�Vf,Z�X��Fc)���G�{�If
U��8�X�&&s��2���S�=��}���{�����z/���w������Tj�JQ�)hfb����`{[K3nt����'�T�V[kW*�x��HcK���ԉ��XX7~��Qח������_��y��|�㜤��λ�N�tcN\�����%�TP��s�&KVKo�^;r��R �йfdz��cj�q[{�T��qN�g�\����ӫD�gfZ6�+T��§�Lv����
�bqS���\�x�J2���/�y�Ď;v�r��?y���6͋��q�J�C��xi�mԾ���+#Sb�nn��\�v�}ͺ��5�nL-�R�-c�Ղ]/�v�s"l�<}N�@(������j�s%����ٕj��C�*V&V�ׯ��FM4���7P��D���_�]��$U���DT��.#�N.��b{���I�o��i��J�<{�Ʈ[��-k�cj|��5M{�}�{��ȭ�*ټdՅ�갾nR�pM0�c���&�y��x�ƹ��6�4�<>���G;֭����qܷ��kbe�1⯿{�Z!��Bّ��l�S2dS1�1.����M6��;z����WF�H"b�9y~������13ٸ{h���ݣ�����so�u4_X�&)��s��OqT�T������
���%�������׫R�0:1��G~��f��O�p��A��H������F��-�JB�Eߦ�,��T*,�:,��c�7س��R�^x坱����&gO]>}����C�k7_��~xX�A$p5p��j��Y?!M<����eƛ�����#Vm/�c?��9�rǁ�;��5������_(qjrr���/����?u���o��Z`r+E��͈�ӶύO�r������Ծv佁mC�ܹ����w_y��G������ͭ�:Ͻ�����/)��}��[�Z��+�z��U,5:6��/ս}}��<ppR�0�}�7����P^k��^��/=�4=��_-��pB:=ԙ�4nd�{�S??z��ؔg&�2|/�d٩�<����V���7��P�^(T+���6Q��]�[�D���G��9}a��ٹ���U�4��D)�> <��+����b�
 ����*�Oy�779���-.X�l��I`\GU��?~���d:�m�f"��_9z�̙�YKO��L?�kWn��3�
7���u�0�ڶ�����4*[Wd�w|���
�z��XD(�qo���B����T�Ȓ��r��W^����~(\`����ohj:{����\��X��7����ᓁ�tU�����P�a��+G���'C��?��lٲ�4M@�J��?=������<��t9��{.�Ӄ�fY+ī�K�П}�Y�y��Q ń�6x_Vb@���s�O��^!����*~�T}���`��Hx���I�����F���_�K,� ��q��9�ƟF�V��*�O7�����Y�	��W�W<��d��}�]��h:K��K}����h��������9��_� =�&�����R%J;< P[ʈP��N�#�Z�dƌ]�zU�S�0$�VHt8'�s��(����a&�� V� &5������w��v����kTZ�gp�dCIW9���A0���T�Ã��������)"�1iV��G�^�t���B���~��uFM�w�\�a�l5�9�lw�`�iDZT)�hT�x��%�=�B+�k_��:=9���|���.dvzkD�,�C�0�${��\�,������/�35�Tݰ�ڛo��+ύ�V���(B�%vV1�Xa\6E�7�k~�w3��c~ ����ڕsg�^EsR�����>0�Z�������3�©�A��t����hN�H`B5X_6:T�^�,"�V���W�z��1�V����ыS9�)�Lb��<�tjfz��3�����&�.��O�.�#��_ʳ��◿�eS%�����O<��/)���%H���q�*�W�*�կ~�J�Ka��j��٠����K@r��{�+)�DO�/�OXzX��3
ς�}lrÃ
\�<�9_^\�G�p�e_���xS�%�N�#��%���SM���"�:�7��/,`!�����k*1Y�I߱
ЗR��FP�.D����~�F/�)56��a��G�\���)���	f�6Bt��a@FF�)u��1�D�i�1�� ��l�_�E�J��<#3&ϥ�EY�2��I�x�����;�[+[�+j:Q;iJZ�5��C]��.�3p}����
$ƁW�X�Zsu#�r�e�a��n_�f�KD}�Ze�����`�|�Ȼ���0%��U-<>j$�/�$b3XJ2��[T�긁�E��� ��v��"P�&��~��0f�|q�������^����&3�);~�j�[:g�
��y�K#cX]Q���R�Q��+�IQ"};wy!g�L�V�3�Ոa��˕�-�XԪ����W(+�−�����͙l��xJ��}ut����������yFD,*D� �Et"(*��JR>�p6qB��ԭ���x�H�N�M
�W睫/T}p�D���r��T)J��N���L�dPp+������ř2=M�]z2��e�W�S��� ��Q�W`d�bX�fb����X�bbƏg�4����]��ߊ�5��g��'#�x$sel��嫪I��]�{5�5ۼ�H�E����m��-��LF(k��U�{��)ϩ���R�S�/���"'h���fMN�,����D���h�3 �
\O��H,�V������-JCP0Ö#Hn$��z}beeeӆAܙ����I?����l��E|T"��9�ٖU@l�g:�(���J��eψh�dey3����X+� ������Q;ԅX"�HM�Rvv�ֳt�z����9;��x�*��5r�|&�H����������t�K?����TA<N�U�2���8�z�+	ը�@]�Fhkf�iA��hŲt�ֽx��*Ϣm�L+,�]� ,}����Q�{Ϯ"ġm.�ĒW
��S.QmV��L��~��{G#b "�nQ�t��3���۝ڎ+��Z���O�ą ��6DVmL��J	S�4�I~��17�F�d;��k����<���Ш�r�Vm��ɯ^���$���D���r��6�ԯb���R�3��3"�z�ѯV�ǧ�d��� HA��K.b�p�ł%�ƬzČ�V󵓧����ߴdY�$_U"j$ze�zqyV%��r*��	�,څ�B��I��DZ[^_tJ��4�V��0I~��%������~�)$��#����}AÍ��l>�����e�419�626Iu�6�R�7�
�g�-3��y�m6C��0���mS?�\>O$��� :S�r�}�xV���̭�ފ�����-*��f&IJ�����W%��P�\���|b����3a�|��C�ܮ������jFMBі�'��`c�O�Ub�Ly�
ipGa%$KaI��b�ؔ���Dc�)��f���e�Z�T�Ny�6����&u�b���X��_��Q�PzY&���*� �Y����M�,�DX:�Tb���h��s�b�N�,=8��d������٠K�]����F~����]<�LLL8�2�N(hS��f����J�&�!b���8;�{w��g�ǹ�ʘ=F����!�'f _��BtB=�8����О��D��Ʉt�ĕ���D���R+�J��
 �%�5���*�ݚ�6!t�~��!���!N_}}}+�������O(b "��}�z
��aq1e�+lE�c���O!�`�b�
����1�0o
�G^�,n�0�R�c�JW�1�.�E�!�g�ԩ�F��L��i1.Bx�(��rph��FF��!^�KC�M��X����p<�)��(�6T���.�
 B����
�)7�6��Ya�E`	��y���+�*ܸq�B��[�����:�	��+�aa�3�ݔʢ�xzn���Dt�G"a���κ0�2Ž��f(+�!���jQL� ,��5�:a�/�"a�,�qٙG��%�F\N� w������l,��3#�Z\ΫPj\n�����7�Be�<�hlH�"�&��̄6&��l��54���^	�t�qe~e͚5�l۶�]�Xe����Cx=���g�i�^��TM�������4P��1�?Σ�_�4E�U)e���I�*�}Ū�m�L%!�x�-�ȕN��S�8���>r�_|������rJ���:KB"� *@տy)��Y�Fu|�JB�Ĩ\��^���Oza^a�0b11.L�ME �:{ĭ����R�}�ɕ�EN�EQ�'���$�IU��:3�������=v�`����|���
��|eeA�M���E+F%<���k���2��פTS�RnX'u����^��I��B���4������A�T���h���2������lcc��+}��%�`��>U3D��r�A���D���6�b��2�<��V�,+��f3S5@̑}[��Dy_)��M��ğj��h+�dht�>�u����1�h�bt|jvծ�K+�ͭ��hD�*�h9����ϰN����3d/S�ڪ��u�p��D��9�af���L�n�B�8��zR�������z�5�|�4�n�Ԭ��	5�&���8���B��[nO�{��zW#"�ѥX����,ޡ�Ź�d��s�e���PbF��w*K�����R=��7fT��G=#�l�Z�$#��,���JM��-lذ���8�ӥ�ׯ_�c����bD�(-[��ߠ�1�`	Ay2"7&���1C{�@@��2��;�b�]�7f��++��¨��?�B}��*׉|"P��JVQ�_�+~=��bx�h���8Ѯ�$+������1K�XX"ç�K��-��
(ƻ��.�/Z�/��M�O��ȶ]KFk0�Z�	Zc6�ˍ�zZQ�*ی�e���[U�PZ	�dM0c� T2b�q�G�+L%Gq��Ng-Q=B;csK��256J;�Nū{�� �����J��NS-��U,qq�	�f�o5��Ѽ��/'�_ϗ;KSY�O��/�)MMX�z��S�#N|�N.Z5^1����S3ш�B �I1���Vcm��2S��r���[��Z���آ��իW'����p�N��c{��˅��C��E�H�m�FD�:�ҠQ|��y�-�B����\A�F�ѸF}�˫S�@�ͩ��LJ��U��<c��|��ϋ)!	��d��*չ����\����_|��v�jJ��jUQb���p7�o��e�+Ǐ�8q���uG�j�2/�.��&���ϑ��1dD ��їf�� � ��R	��Q���r��nܸi�Ɵ���'�|����yOO�e���X�2=�CC�Y�k;��6R+ݶ�N x�l�(LG�r�����<\���� 
p�c���9#2Pr��93��ٽ	/~��A�*��yޜ�1v��) 5|&l|�腂0���qxdܷ���:���q�w<��B�?n��;��IO�s�:�^��� �H
*���� r��)�<���X��L�C��&���Z2P�4;Bȗ���.\�|���Lc�C�a�M�e���'�YWv�NF<�H��ر��!���hY�T��Çw�Ǐ�e��aJU�)��I�!)a2�K䨳.f;�W�L1�Binn�c�F����kG�)�"����m��lVh,ܗd�~s���C������IR�ܾ�ۈ7�Z;v�س?�= ��Ӌ�^�ˋ�]԰�$d�ƍW�]�ج:�{~#���	��jn����E��R���gO�>���^�q�02��0-�m��$2aްڼ���bX&8�Ƅ�s�N���_SS��Ʃ���p���� 9�Nׄ�`�1��A��1}��0utG�������L{{{�z�����*������9E�R����ͭ�g3a;���p�G�Xl��V+���w����d�k]�(n;{ys�s�T��7�	����iVH�ʳ�����t�,+�ցu����-� ��5��g_{�k��+b2UY�s>l�g�q�s�7o��J�q��A�wo^�����R�
�K���N5�SS3###�_÷z���hQA�r��+V]Pmo���땉�������������6�R����k��4��s?{sfff��v�*	jU���WeՆAxDA����$uʸ�ZS ʚ�~��z$�Q��F��;�^�r���]�H�n��F�����j�H�d|~ϖ-��Ƿvu�`���=��>d��lm��={�|�'/b�X����ʿ&�������Q.��`��v�e�j�u�Yڠk�M2+W�1s��5͍�5�s�EI�%H�j�Wh��;v����_����T-C�F$5� )"�I�>T�АMۥ|17�֒^�nͽ��P�� ՌFښ3��Ļy��ߵE�=��0�YVp5�sX)ևѫ��0��c#X���Z���
+���t�_�n��}��{�>�싯�T))FS�Ȋ%*7�m��x�U���J�l�-c�x�48@"���Dbjq�͏=|it�_��_C����È���=J�Ԉjey^��j*)�c|ٶ�8��[��8��YF����ڬ�N3*��܍��e]���ؕ9�戼x��#��	�*|��Y�n'�������7����#�ǣ�����c��Q��6��LOOdۻbFd�*��#
��ϷeEQe���
p��%dAa��L�k���m]Ӓ�"�&�L�LMc�[wm����_E ��BY�y��Ǥ�����oa' h>� ��,����d���!Ut�o\S$�nPB�������z뭧�w�%�NzdC{,����ʙ�{c���v�/FT�S��R�w�ĺ�2a<�G#������������Q o���hS��HT�����m��h�Fs:J�8��ys?�L��W��Hqe�9kg�E��lNE�}��o����QQ�]O��z'�ATyQv����Ej5_�+����]�o9x;�F�^����3�>x���я~t��o�-�1�<���7�>S\���B���J<���M��(��z#�I)�I�~�1ٿm��}��>v���x��^�G͈m��h�����Rf-!ƌ�n�o���m\���DIüG'F�9�r���O<��E$�ljr���Q� �
�z�m}n�Fkm���rw����w��APokNu6H�Doooؾ}`���SO=UY���U3����ĴoբZn�V.P%�h�N�	�T�/�hm���}ǆ� ��h����1��=���={w��=��/�x<�bi��,��΄�8� �d�\�g32W+W�vu���s�6 ����n���$$)]�������ԕ������H�Y�%&��[��dD���]t�zM��==�x��m�k��昑'�H��`A|���E%�~���\O�X�cy�ʹ�o2��Cε�%�<;̊�����c��h��.��_(o:BYw�ĭ[���o�ַ��-x?�w�N(g�#T~3#ȷ ���P��n�o�-O��)t\�Q�k�L��}��-�ܢ%�_z���'.(�MU���P!"T궓��z��C��ݳ#��gѹ��K&��=�(mg�<�H0�,���D�R���
�ѕ+�������|x߮����8�R�R�9J�ضm���w~�5�J�@��>��:|	̑�M\a�`?Dy��~���$�j�f��5a9������k@a4�\(��Fqޯ�^���N�d8��!M�k\�Z���Ij2|�uy��)c��Gҝ�������N�O�>��U�{����F��f4J}wKej{)h��m)#%����z�p����~jEݾ��ʘ���=�m۶�a�
�_ �6��2�Wزe]6�͕|k�U������?|v:%��0�)�$�g��ߏ��ˤ�Q�j)���h�X��������5�駟�=�z*IF���6����'��0��n�
��9�&^�5QU���������X������\N@YmGgB�|!$��!R�n*ف�G�B&�(��a�:J2!;Χ0Y6���/��#ufU�z$B8����a1>��oM15Ԋ�����5���8��bIjl�+Q�����B��_Q�XS���b�,�_Ux�ӘN�
�-ԋ8 ,�M:JQ�����,_��~��<���,Q���sT�7Ń�"-x�#�>�я��T4��餐hl�B�y���׾�$���)��D�ű صY�
����8?�߷o��J�˾�|�l#�3�X�"�R�s��V5:1
-��tY׍hTϔd�Źih����x mR�^���y3�6Eo���[�{�L��딉���I�6&a\�nb~�S��6�Y�;�g��vɠ��������P�̏��ݺ�sg�9�+`A��Q��`?� ���[���`r^%*h�1�=x^mv5� n]O/�J��/�&�V��5('4kH�p�j��C{μ����vU�NCUJ�ǜ(_,R��4;�`۶mx`�V���JgG{s#q#k��ݚv}.�[�]�~ٿs����W��h����tꫩ���G�:� 6Wen鑇�Ø�q��Պ��%!�-���汉	���ޜ��O}b�o�N��\�<�EBl*����p�EXC��e��y��W���;b��[�Nʦ�=�A�����*��Xa�ڻupa9����[�դ�M/�r.%K�@q���%���:Zc�����x�ݻb��0{	*שi�fRbAѲ˖G&�ч��~qve�T���;������|�)�H�K�[�Dӏ�}`c_S��
��jk�zc�͍=TWV[ں�U�g�׾�D�4�>|Ę�!j A�j�_�^�zq٫UzZ�l߰kpmVH5M= �v3���K�J~�Fw�����W]�Eܹ����V��E��Tڨ#Lp����7x��&X�̶�X�����Y���3������|R�?�ɏ�.L^�^!�V��E3%TjUIQ<;5����_�q�Н���`~<cJ�l6�wT��<�T
��ܩ���n(�����W�PlO0�f�6�i��`�i��y��Jp{;7�kM�����4aV3	:9��ȝ�u_�����^��|���JW]'��K�x/p�*q�*��{�Xk�Z�ܳ�����M�1CoiJ����v����b�r������0~�!-Qo^�GЗ�e�D#tl^_������w.,���}1��"�x�R5{Z�r�23�<9?2��5����_���Ja9՗V)m�5��4A�#U5�Q�m#jmY���!�ᢲL�'&m�񈙌5M� �&&'<t���
����>u��\2�2C�Aū-W������-�U�^�Mmވ8 ���PQX�p.�R@]��xp�F���/}�K����dģ|�HEY�U��4��@m��ܱoS6ʩB5�R�)SS�:�@����������~�����o_M��l�ui�^�چ�r�\�lY"������a�!�u_ߖ���O5(�8\�B�S�k�������m��f�O�_���Tek�"����Z��B����V�[-�\�g�S�$I?�l�����C.��φ1+(�/�*�m���]).���V)�F9|>D��������m��s] L|4l�~�0��a>jPu�޽{'�t�C�.u��s�-����R)���o�W���6��V�Ɔi"�(	�l
X���{��+�υ=� >�L԰�q8�ЇDp�/�,� �B�׭[g5l�H�҃�Y��3�[�Z�C!uj���V2,49d�5}d����f<����8p�^Y����hj���w�_$����ʍ9,��呓��Tn��� YЀ��azzz�z����bT�������#n�rJ�ڪ"2m����ï߹�z ��6�
;(���$�u�"#'O�q<>���tKc*d�ST+�_/�z2��4��T��g�X=��5��3�%������Gc�(.omLyB}�	�F"F�v(u}�PA��|a��ɓ����
5���!�g���� p��l�C=D|�	(W���!I��:����=_�`��l�#�<r��E�_�Xx�1�!ک����LC��u����/]&J��z|�̹�bxv�g���KW���"$�������G�	{�sL��6϶q+=m�j�7��jX�t�R$�(�RI$��T��^��X�Ls�I�9��C5��F9<1b�ٶo�ؘ,+�i<��˴�ӳ�0�����Uy�ڵM5����P��}�c���ˤl�7l�� �
��� �-q-,XٴiT8�j�o����twG��ק��� �N�����橗Y�y83UR�y�۰a��������Q��Ws�XL��(8�?�Rb� <�UY���gy�,]*����vd{�1,(�={�Pm�L�*Q´�x�qu��ǎ]E@s�=�^}�����{����e�%���F�n�jm&�ggE�f""���9�j���~*
eX�2b�>��ϟ���)iXkB�3A�� ô@Glƈu�m�A�3�,���ĳi�"�+	ץi�X��?>U@���W�tͰ]�i�����{���T�!0e�n}x&(!O����>,��<���ޔ�"��tU\:R�Wr��/����wNd�W��!�|gby.�?��,PVA@��|(�U�۞��a5i�ad�
���7�zgz:_��t�E�%QR��ˉ�\���F�zv�_33|��9�֔f�B܈*p�R���JɳqE�̱�����u�m�.��xc�fSB;��d٨5��F�����3	(�Ɓ�Z��Z�������Z�FS�L�Wi�hpp���k��mS>7�I��H�7g早I�tC���~�^�HA& k�G~5��7)��c�6OL�s�=�6_���~M�g�I�(`�H&)��Ja�Ё}����]������8*�N��K;�rS:Q�ղ�k[����ٳ7|!�vx<�y�3�¬W���=}�]{T��?��h�ʹu\�F��V�����D3�PT]t���m�N�v(Iݮ��%ip{��X:��[ƈD��u�wh�Z۶�WM�s�uI�)����*�D�R����[v�2����41�&
�s"��},4!�pK��}pۺ��O��{(k^�-���o�*�M)�QU�h�O,�Î�ز�رc�H�J�
#y�s��Q,���ٱ�rߖ��ƴd�'й�&�,A������Od���?r�����YBDt����@d���m�<\-M�L����rNGC{�>;�"Z z@�N�V�{=�I��/~qimۖ���{��iC��"ֈ�`!b��hl�W܆læ����Lc�
y`aKs+$�	N-"pZTK�����z���p.���?��P����@��&#�nO����ե`nH
t�[��,G�ބÝ㫜_}��;Ϟ8��-�g�VJ	G(�N#�p��j��}=홖,SĐ�[�9	���F�F��U�u5��93���u���~��0���*�8��D����9�)Gx��!���9��W�W	���n��۲��ѣ�W���|����I��P�*��oB�<��MD �K��P���ܚ�i�gJ���*�N!������ba�-�n�oy��À{�6�8q���t~)h�իvT3x�J�1�\����g熵�/\�(i)�r��P1���m���u,?+|�c����ϗ'��y^xO%X��AM��i�l_�ɹ����|�(���j��+A4�#�H��=��-}s2���/y����~�������(������y�	"{Rd������2��0�+���a�+��j�933��<���n���|>�q�F��)[�BX�M��Pm��%���E�/�@��S���cuC��?C0�H%�1�i�8�Y����k5M�X��j��#˗�F���<��1x�H� 0=��e�t� ��&x|����ޑN��m׊�]��]",O�u��Ihpw��c2Lᬆ��l�_b�թ�)��\��yq�B^c:�Y�,���xnu�����@K�"�f�\s�l̏o��su��w,^4`��t%`6N��pQ�M����0:1�I�Q^A������
E�"�30�Gt�����R�:ڽ%4�hOJ�Gkcn��n]�G>����kk�:�0%7�pR��E�v���l��"����/�B�v ye�����Ç}VOı��:��S]����{�n����]�U�o�إ�6&-�a�����Z�]�QE�/�����y�� ��Hx��"0�r�0^�Pt��3�m�P��[�eD3�;N\���9g{�.�n�ϫ���ԄG3Mj߆ϨI C���B�űH�4@S�����bBz0��:�He2 ���O�,��wk�ZRV$�"α�]�f�	:��-���)�_���'�\aHU-��y*E��sN�5"���zE�^G"�R)L��Ѹ���8������fc��JdC6�͉�X7�I�0��Q���K�	�9����^��d2��r��m�zble̲�(U���tzQ,"B�г�9���ʐm�*�is���wb��ؐL���\YKK�¹��S�GM`�?Ԙ�#���q`���l�S�oq�"�3F��?�>6<M���M6��T0���L&�12��z��Q!1�&ߵ����=p��RQ�B]�0�"U������I�������]_Ue]UK�Q��[L�E�ZIS��C��Xr�^�^������$��[�jk���,�Тl6{��Uߦg�-�A���*V.�NȬY���-puMf�.�-�ܾ/ҍl�j���3u�B��C���M|���(�d�僙�Y���Ri�kk�5�*�~ӧ2ެbQMUR��MΏ/T�ħ�P;^�|�ܰ�����K����b)���(�P$��I)��kI�QI������̩c�,���fWKrܤP��%��I7MM�dt�lѪ[*�S����0R�e(	��l<�RIה%V!�Ǣx:�nL�U]TtU���Ǻ�55�����D.�L_$�L�mjJ�lE#�bɛ�|Q�J���ձZ�h�T�U�O�m��D;���hk�$�ɨX�4d��\_��,�h��JҾޘ�͏tQ�FR�3�y�*Em*U�Z�]�R-7�Q��nmjN/-�54�x%��T�;�\/�t��-vJB��)��RJ<j���\.FS��]�4��y����ٓ��x E�T����^�*e5I��\ߓ#D˫ ���fLشy��<G����|2�Tv�$��]5A�����İFMi]ڗ��.��a貄���j�ٛ/��o|æ/^�i��#�X�,תS�Z�Zm$�1M���V,�_���)�KQ��p�J� nU*j�t_o���y�֗��� M$�δ�����Y��ޮ��ˮ�R��N�
\�
���Zu�2���9I�����pNsK���uU�<��[C�h!�F܄ᳪ�XOZ� �6��wy_��)�a+��D�UW2��}k>�ط~��b�,�m��zHV��N5���8)�DM�(��)��O��m����#j���kh��-��^���4�F�f	��L�G^�T���|��dウ:%MpT^�X��-�u�dS�D:���4�&��;���g\u��`�1@,yk�3#zZ�OO�X�������y`�pR�yb���T���dlvr����|��J<�>�B�ZF8�{�d":?s�)�RU����-QU)֥�fV���T�)	.퓱�5��E[�9���:Q����^0����nt~BD^�wCtV�,�B�F�μH�ڗub/�KQ-
K'Qf۲a���v�������H��_߇b>9Qk5'<�ը!�����2~�p��a��2�L�k<w��ݬN��HI����P�([1:P�#�Ŵ��F��(��$��-�D�����۶7'�N�Z"����z��&���4V�p��5���Of:��uj`�cr��Y�:�Lm���I�d(>QY�=m.�!��ѺnM��Jr8�Q�_�����r���[V�rIF�V%È�XM(�
�9<N��1;��dH�*Ўj���hNY��K"��cM}:g�j��R�N&�aRǶ_k���Y(2w27M�8���d6����j�zoQ� �>P����𬼜�3��l��9H,ڣ`�H��&%/�r9���q[��q��ݝいUVa��F��f(lT�g����+lf[+���������c�Ar�ԩRT
��Dp ?>11AP��]ͧ1!�2������Q�@��ݖ�V+�fF͛́C|�ۖ�2@1(�#�Ά�2�n���ދŰ�w|||� �O��6�dշ�i�=������ܰ7,jA,�����1r]�yoߪ����6��T��H��D��fg�F��4�	��=@� � �� �G ���dq0�;��X3�m�]�Hqw����fwWw�^���/�;�������,�k�U��w��|��s�]؋>\`�
Mް4ɄdU_���cN���L�"��6�h����q�̗�
'g���շ��U��L��F��A���'���H��v�`���;���N���2Y��pt��Kߙطo�R�#�!�� * ����Ge�Ҫ�U#G��F3��!�<��$6Q���s�V`���͛7�5A�e��ևGph�i��s�( v�-T�*��_r�t��{�'�� ���
�]���F���PS�(��I���s�-���Mh��l�(b�<>"��/���H���ЧQ!�ߣ{�Jk��^/�"��v�H���^^�6ճ�=%�����%�Rm��4,���-�/�i�͎K��+�_0���GJ-���;��z1���{����� �A��K�3G�tʇ�(�W��J������ܱ#�v���D����<� Y����l���4�	`H����a�pM�?%�R��5�����X/m��F�r|Y�Z��Ihl��诞����$��S�Oz�c�8�����g�^=���|�mG��HqD���L��#<q�"�;7��d-55�o'�Bm������9U7�3�7\�Y�斶Z��r�(r��=T�	S���d3ق��ӆ�:	�CHuD���Q,kV��'�٩���b��^�����G�p
��vA�iغ�1�\��V��UEs�!�Jb����F�$e�>Ti���UZx��i��a�I�O�d�3Z¦^�V%��_�](a>U���Mryz�X�ՎT,�F�s�T����/�0䘆�wDf�iu@MO���4���'�,z���K��w�j�2�^@��� `�,�Zm������d�'����`�V�m��@M��4u��U;�Pr�P��N�&���\vi`�i�n�&����@�d�w�\@Ɖ �ؐ��������뇎-ӳ�7>��ъ��K��I��m���ZmpW6F�N,G��~�姻$��(��w:���#_8>4j��z-;0:hYs�Z�'.��J������n�D��*�K�G1y��e��d�:��z��3�z�����PR馩���1	i�"�N�+nE�-Z�����3R����2!9��ɡ��a.zK��@�����e?���;Ȇ�5'C���̩K�c��6���/޷{Ϙ�p��HK�$��=P�y�����I�Lͮܘ�&�~{y+��٦;��:RK��"�.	�	{�;J�Lr14<�`�m)ۜcJ��2Nt#S�]��ҭ7ʍLnPճLi��ΨO�T��J��:ع�[Fh�#Q���d�a�U&��D\F�ı��+�M�E�V+�<�Z�_A��u'@bJ8I��!��L�7)�q?�ww�F]%%P����z�`Nl�(��jm�7�x���={�ɖ��oIr�|O��nJ8�!�DЭ���"q�)��Y�6���~:��c8"{����M#���� \.��B$f�"U��i�Z��2i7oU�ѥ*�:��W��B�m�6��n��6gkx���^���{ ![E�%�U��E4����,R_n߾}��3gΐ0�ϐ�����4�HI!������֦�B3Q���SB5�i	bE�'qHCs�^C��������=�r;�Ld�6��R֚��4�3�p��E�	���ܹs_���h�/_n?����"�k��(d(,�ѥҖa�3	�c��|�\-��+)rcD�ɏ?��T�h�� �B~.Hp�NG0�p!�D.���)a��c���"I����E��"�H3�����qCД%�E]|���Yȃ����,�{ފ�R$�F������O�7N�:>�'\}Rsh0Ƞ/�������]�t�8q�֭)�y{�8���f��b��״�$~4��>���c�H�ԛu�̂��M�x1��pnii	�P:MN5�A�`��j�肴�.^���K/M]?CHv��"��IXR���G��$J�-I��2|�N�s����/*�u`)����ٳg�?�E^�,�;�k+�1lJ�}o0�޽{�}�]�{�F(v=>]MKz����ȕ�7r���L�A['E� ���ћ����Ͼ��U����>ow<<�N����U[�~�7���h+.-�Ѐ��@�Ռ���_�1368z�E���열s��ד��k�:a�ѸJ �'Dπ���>��-��؊����h�5�U��o~���O>�D�'K����SD����fU�3�D!�*l�X��9g	�o���J��&�O���9b�;>�@�
W����p���/U�{oh��X���0�>�yc|bL5�v�M�qb�ٸ���@ZY��>y�l9U�ݪU;�:�[������|x�8>����S�N�oVѮ=�&w��5�1q(�.,l�ڤgK�F��:s���$rg�����)*��{'O~�}C�f�n�يd���N���8F���Nim��KwV�ݵ�����c��(�1dd��_�ڊ@)q��y���=p{�О��j��9DTR�l���s����;���\r!c��]W���:��۳����^�v�[_��" M5i�P�R�پ����[�&zń�uG�)�CZ9�@���[U���������W�<����xՄ�K�K���.-�-/�m��oV+wK��D b��hUM�<��$�|�T�u��^[z橁]css7GƇv�A���4)%�7U1�x�:�Ų���l�P�q�i��dr��8%R�c�aC�_���_|�藾���o���of�V�#��HG���2[������}6�������<�UH�e�|��g��T`�[�_,o>��7�y��|d��$���G.�A�8cpBb��ҥkWn�>��Cg/_�]ZV2��͐5�Dխ$	�}	� ���������WV�^�z��\��^j�L���9��n֚7���(~���?���U��J��#+Hv���гl��F37;͙�ʓ{���yet�xqh7�k�_	8t��WZ����zeqm��W���T�:�`����{e"ܧ7%�,'n�lU��~�U���s�}��l���}�Vo�*�]���n^��x�Ň}��|�}���F~�f*(.�Bp�E������/=q��{�&�A�E�C�i6]'��QBJ��g/<����\��Ot˗�0aw��,h�+����)Z�TU;C��ܧW|������,�$��x��z������������ݕ"�|7����K��v;�D��0X�lV�fm0šqrr�>Ҧ$U9����S_��3�����z��9*�ݤ���h\V�����Դk;ٍ�fi�������N���4�i9]7t��L���O.HF���}�|0u��Q�ǹ�!����oEA�^%���7�<�_UT2	��E�(/�,��"�[fDID� �2,��n,-n����Jj8�o�U��=Ug�?l�]R�U2�QaY�&���w(cg����i�s�+��&cH׮][XX�ߒ�%�	�9Fp":Iן��A��ONN
<۽���f�@q�T% ?11177G�4��ʌē{"��4��& C����Sǎ�\�&�:��m��Ok�81_]�_�1�%�!�Ƹ�XFD�1��=*J���8���w�96A'3:>^/א}i�J3�g�'O�����u��������U���!��0��^��˗/���s�}�.�YLU�z���Zi��H��خ'N޺uK\Mtz"�����H�i��p߮�{�ҹӄ���+�
B��i�5=���X�C��H؍9 �'��Т�� J�i&O�<��3�(�M�-�Q�k1Ӌe�����;w���:tn�.aCE�~��Y�LA_��v�r����~�k_��O~B�p��фQ�c;�tm���3�$]��^b�8���5N�|-M(ŉT����5p�|�|������A%[��++�SSS�?B����oп�8\�B~��{��nM˴��������Q̪�#��C���[$$�"�;�9uc�V��uNe*Z2��K�a���%����!��0V�o����"?�|��>?��M���]#�gN�찘%R�|�� ��qr��'4����4����B���]����F�s����?��ɧ�AW����&kb��F�b����Rd�DO�|h|�FB.���Rlgv:��+��$H��]���ׯ�Qԙ8CR�ɬ$>�A._��.\ ?�������q�JV�&Sj4ݛ7o�׾����/�~��_
��nNH��EUm� $��B�J��D��S)�=p�����2q�_��+��z�-�~O��\�/���@������4=�����#��O
mx�(�|9�Z�т��{�ѿ~���R~pj�p�V�:�:!��������o�]G_պ�\A��Xb�	a	� ŸѨ�����n��|�j������G�*��!�[7��p�˛��=4��(�R��/\��
m ��a�6�w��l��_(y��_i���I���8�3�i�y+4U�	+��٫�Fv���ƚ��X�ᤑ���u�������y*X�В�H�HeU��c֨�Z/ �p��rx��ܯ��Q%8s�v�7P����8�ܘ�:�G�& |�-�C���9[ k�r6È�j�����^x�K_����</�T��jL>�aC	�}`uc�����'���|a!C-EBs%!&դr�2ؿ���~`���Dsk�ެ�-$��z�r�%�@K���-/m]��Y�[����i%rL8s�X5���#�c��ʻ'�����74>\�mȊG
%J���s�|�6y�gr��N��xza��ZVF] �hP�!Gi�˚��r�y�̅��v�G5YȾ�J8ڨ�kln��@����j|r����R� �t
�M9�/3	h;���������o�81��|�_�l�K[u[�8�Iiu�Z�B�����?|ij�W���y�{��`�U��E���k���FZ�d������3'���oߺz��K����]�-/�nllL��!3�{�W^�p��kGAَ38"q��M�ʅaF����3�vOo_�Za�)/ �8�%]p��*ً�1?���O|�Q���i�WJ%gN'�rt��{$����O籃t��h���q�-���^ U"ٹ=����S�.Ǧu�Z�Ԝ�6mJrU5E�<�lg`q�����O�_�������+?��o}�[�'��rC��Bޮ�ӿ{�Ù���Gx��?��n�-�����k�U'C��h��㊔Ȇ�;��j�����t���o��}�>r4h���y]G#�7��/~�l�[�~�h{I���4�'Lގ�Cʹ����H3|r����Dq$����m_Q�谲^"]k��^��3�,����߼���V=Tk6C�qn�dBgB�Z�ݒ;5����k��_y��#v_f�t�0D�/�h��y��i2	�C_z�ŵ�������"�^r*�����>�@�vB�ҍTR#ҥ+��?������ڵť�ɶ�o�>v�5������S���?��Ϯ|6�W�q��m��#0c2���15�w.O�z�����	9�|d�Q��w�i��u��ڨ^�Y�[)/o4�\h�4��ת�R�`ٖM�dY��D̄N:�0�,��5�����߶#I����?�!�|B�w���!��P��3x�A�ҥK������� D�ZV+��ݻ����믓y$��At���1�c�8�G�X�"���D�x�_FP���X�df|��rW����?�яʕ��Q�T��������`������:�ĉ�R��SO�����"�-U* wIHHG���JN��&5�\G�Œ�=).!sS��׿�5�Ľ{��5�8�����$�r��+������C#�|���W0�V�@g��&g8tM§4���J���1�NJ���iZ[�Hd?�p�?���7HWpCn���&�fm��L��eFL4����s�٬m�h���7�����|����Z�{�w�~�m2����\�P���xܺ����t��ƍv~��~��Ps�o��aUE�f?����/p��#��qW �@�T�mC�8h"Z}����.}�������\�!]�[�ڦ�{�h~���7	������HLZ��zK����v�|«_�{�s�������wFFFh��Rd�ס�1�̳�>�������++�/"G�}1�x��L��j�C[8Q\����!�k��CIۄv��"I��UFb~��ja������kt��Z0��Ւ��Idx�������W������O�:5;�Xt�ϯ�YE,�?�x��cZ�={&��D���i'FX�9�MEA��uE�+��7� �r�
|r�]3T�nl�������_\,��~���ؔ3|�8G�H��e��j"'���������?���{z����L�͓Ď��%�-���?��!�� �4;����B>k��Cj�������W��}��GΟ!���ޯT�4���=A����_� �C�,c� Uk@]�J	��}�,��/��/����d�V�D��O�ܳ&N�=�$�������/{Q�y����5�nG>��nA�Fc�����#d�	�*��sd�td2�����M�&�k������ǜۣs���#M�UIu��D�����ުk�;��N��>��i�M�(U7�=�(�~�fg���J���]�N�����_�[������h���Aa��k�5��άl�����vyy����㊔5�ut4����͓�_&�7u{)-ɴ5	|�t�;��V�x=A�&���[���B;���^Z���0>�E�h���.�����ק֚��4N}@Zd�e���e�
��ə�����rN��i�/��l��>��#��A;#������W��9����\9�Hƍ�M˫Ţ.��p1�r��Aڻ�4$���\��ڇ�=�rr�?먦�GRa�ܒ�f�=�))�)7��޿J����{���BIR�0�p	2i9I���H��wO�,mŏ>�����佗���(c���������]�Z��ŹB�,�Qncb%�ג�2fX�k���]���Q}�������w
� �ˡ�~��S�Ή��?��/I���dL��}d��r��s�i����,YQ��4k�F/�㕗�y���=*����V��9��3ΠZ*��:s�^��� �&W/�K�  K�fxQ��n�W��7tZ��� ����+[�~���}�!2�n�/���``}��x���oܜVr�A'M���bv��L
��Qd�Gٮ�ڎ�uI^�S.��k>��#G'���n�-�h
r��)I}��ۧ?����1-%��*I�R��o)ֳJ[8��ݞ��H^�޹R��)<�H�D5���g�w��O�?YX8��I4�L��t�\��� �����ˤh6b5Vr�V��c�ʭǪ��q��8pt�.7�pRiJ��S_��������edt��%U����AL�0f���6j	��MY�i�YI�]��۔~��FJ(��r%�9�cǎd��oN�x���$ݵg)�|� >!�k�e)���y�M�d�$$��F=���9G���#ӑ�%�ˡ����<F�{�������A��06뾞)JI+���f��w%�E3��ǉ��4��ȫ��7/�ZhI_}�أ�<���@"C�p� ڧ����>�_Uu(����QV53Bܔ@���R�R��Z.�̙?�&������W�z�'#��=�Y(�l��^+�������}���W��r�P�(��غ�~G5���	�m��W���N�����đ��M�ǘ_�Ő4�jحv<??���*����tik.5U/��T�-�~8��6��:U�����dl67�'W�R���#���o�k6;;���3W�^���Lw����D g\N��2¬�-=qb��v��>�b3S�z�A��&��!*[h���I˪�3h����l�������3�����8-�f�E�bi��F�>B+Iڅ�;�=TE�^�r�-�r���^�p������� ҍ�����A|u���*8�Wu�ɓcVs"ACL�c$�l�-6d0�j����0�pY�	��F��Vld{�\����vBm;�."�m#�jbl�F;0P�+���#��奥�X�1��c'ߛ>:gb0Y�C�OV��ل��AҺ�}�ΡC��|�mg�5�,��t�
?�&#��>����#lۇB Fm��Vess�QY�Q�����3Aҵ�Q�}��ti���7Lf)�9�饶HX��b�-8������1���&�Tx��M��{�z�0��ږ�Eu�� �D��V�$���$B���,�O�$�<��a2$[�kt��ˋ���"�q;�[���v�L���h���VT6�g������A~���n�˛5��0X��c��c�uoN������[u��v�=&�49rf�ޅi
6S��^�p���^���w>���I����w5\(��b�Cpuj�=�*c�DC�X\*�­�=�Tf�=�PQAC��:}��g�w!�ݍI���M�SԌ"I ���H*{Q�v"g�a�y�rbNL`��wq�y�˳SdT�v���][��N�����/�D�ݪj����ĜĢAi��^-��@VC�}���䦐�|�A.Vh��Rxmq��ي4��r�0���%�(<�U�8WGe��0}������������$$�ܛ�g[��ŧnޤ�GfF����o��Ma=b����� �I��V��;�4k��#�c��O�"U�͍;��J(.(@X�*Uںm��Nl�C7��*�KZmt���u �w28���I�%B�X���߽���G�`�D�@��dی�c,G)�	 O@�+l ��U%�]6☿��o�n�qw~u�D�>�yB��*a	�$�/U�����Ꮂ
灤4�$����HLˍ��J%�ڲ��J	�YKV�ST[3s�b�t� g�D#�ϹH�ب��|��yend��~X_�Ҷj�������a��X�b�e1��*1���Dp̀� �w�k���W$��\l���7C]SG�q��r����K��H1b�"���+�PE�>�3a�WY#��j�K���R|���g�iC�\�������YKC2L&��"-�����W�bJ��ҽ|n�i�z*����r�:Y4R��"��J3�fC�l���v���Ők�qN�7*�'U�쇈&:��(ȓ���Օ��s+�\P�^�f)%�14��	���0
U3�ꏣ����B��;����smy��������(t}#�\/da��RD-���k;�A�8GH�$U����J�6��;�8����c_�R]��+z�~�2���q S���Q�����?��A���)�l�.��Q%�Ζ%s�U )F���q��ԉ(�1�j�1z�WF8V�}0�J[j���Ri�V�j���lҚ�`���V_GR(Ј�l_�!_XX��9<TNHMTv�����$Ew���U�ڋ���3���p �Dj����hX�m��;r��l^b��b�mWւ�@+iNW[��O�7�E�I�3a��҇'d�n�t�ȉ�b��TD�m�Ek�."�e�����?��#��0�>'YĲ.�&�RAN-���5X?M�ri��s�b?�3�te9h A�,�Jfu��-�:�?��v��?4���/.�����8R�����Pou�dX�w`^L+W5��Y�d�v�drv��8O�4>Y�Z��{�V��"�֨o��B1��c�þ"Ǩ�T5��HE&	���!gL#�6�,�,�1r�t\Mَ�I���GT�r�)N|�RE�����+3� �f�NM�I�b}�����Â����qS�D��+׫i!ܚH0�'�V�ؖ�.`�*��z��}����g�1b����#�D�+u�$_<a�'6{�OSDm��N��C!r�VA:�s�G �/��jj0.�\#A5��	����8A�!�(J��8��r]���\!ar�x��M�y G�6�
��@J>�y����:j��H���-�Y=f�LэMRS]�~�3�p�y�n#!()z^�$g�Ȇ
�cn�np�e���T79�����Ie'�'�S� f�#�����d!�F�l��Ƅє̐tO���7&��0PL���Uӈ&ݲ�������d,���W��Ԟ�J��W�!�P^lc�n�����HA��Ļ�ۚF�g��~mB�����)���Д泧,���S3Y�U�r�㑸Y��-?��,"��M59"3�;]ا�1�A��0fh�j;{�۲F����y$q+4Xh��#�P�iHP����j�!��X,���	�;<�Td*���H�c�х�h �B��rr8��pF��q���D9�y[0'.w)�� ��E+rT��~���Z�J���UX��1h&�$���II����c�d@���/ݔ�x��G�����L	�]����I�
r�lj���K{&T#��������A��4*�,JFF`��r}���Od7ؖn��a�ފ�9�HKdA��2F����
�C"�bk��\f����%���9ѷ\�|��U|o�2"F��c�P���ژ�#ga�\��F�+s�,p	�Hc���xT����~�Un	�	�UEV�2�M�bH�Z�f\�����8�����'
��H�)�=L�5��G�.V�*).Y�G�8�]lZ6�dp�-{" #�(1��VCt��*qw��q��Ȉ}U *&����%�|U�i
e0�!G����O�I�@hș�hz	*U6d�[~ڔ:�E�~����Rl�7Dc��3�.��'"��w�� ���ҐNN:!��-B���P򲳤�뛛��0:iF��^�;�"AY�u�2��f�Ⱥ�.#νip�B��D�R���7t�6�H�Z]������A���)<�.�r��g��Kc��E�W�2s���
H�|i�����y1:_��ĭ@�GOQJ��B!��k�2�!-g�	B~�qT��;d0QY���4��G���&(�G!?���F#>��)���#/����C$�>P�fs5��+��@�w~0�GP��8�
+Rh5���\@H>�	��C�x3�7����/�{`a2G,�>�d�p[��6'hl�VK8e<�?���xh�d((�#��h^�ͳ������X��
���!/A��*5�#����N�x�8�v�8J��nU��d�Z�bn�.�2�����!0�F���f������ȁ��0��H�T-2w���AR���(�]���EIn
<M��%	P��p/|,SgB�܅��u�J�3�hS�Hx@��������ݎ����ܡ"'ų�iK冋)'���4�#��ܸt'N�ۮ��X�9�)�Al'���J�.�jb�='F=��l���OD���������0�3b�\w����b� ��6S?h�^�?��ߡ�ݒ�����k|����;ˮ	�NEA�}������WN؜вp��?r�ElZ����Ww�J�vij�U���PX�+�LS�C�c��qH�^�+��{��AB$Mt��'�<�^�u�u��h�s��;ak��A�@j�L�0u�H��A0դ��!h����	x�n�E�B]9�Z?��GF����W������]G��3Z����p?���2�b͵ď�����V��R�;��ș$%��M�7�e�'�D��.Z�S�Ry������.��8��C_����*A��#	�w�γiQҮ	��>D����2׬�2�B���$I_v@�J��؟i�<L̆­`6T�,��a��0�I��f�%j��rG��t��ؤ�%3@J�FI�+E�;�$�ǥ�W�-W$E��}SO��j -�l{�}������Z'�I��}���l���D�-��\Q1<<L�@5�ZܿO�)i���@�N�O�aY'��Q�$�q��7K�f���%2�}`��}2�*��s��A֑a����R<S$ �j��5�� ���)�)��p�b��A�DV�3�D�� ��:~Ȕv�T��$/*e2�n1S%����`;�*H,I������,/36y��0$�"��}���s!�H�;p�T�X�:m��(�d�Dڴ�c�5ʠ�PyW3�z<ASW��,��\��5E�i1�T�D�L!�g�CZ/�ѼŒ#��d�a�\d�HI�ݴQ�T�A0Y)���ĉ��aꠝ@��cl�#uqM��S�	�׃|7po���4�b/�T�	-�M�Rq��.�4m4S�6WyW$!����.����W"b��~���;�{r�P$efL+�1�[ȫ0OR跼869�kb�e��^���H�?�v�U5�P��ƚ��-%���f�<������V(��+�.ٶ�Ot]����#�yl"�#R�^�#�et�C�N����D�3r%��Z��������^���YfE�؅���|A��t��"�����M�/7ȍ��>4i��i)r.��W��U�duNU����0�,����0�T��ӧs�*W�Qa�bU�؉|[�����V���5BV�;}����JKJ��m�ɸ^�@��n.�@G\Z�m�yG'*��( �'���$yQT��@)����yO�l�L5!�V�p�*ЮT�8	mˡ}�Xl�H�J$�=)b�12�>��l��&��;��q�A���b���c�;a�f4S5t*up';44TCWz����:��X�P��1���-G^�f��aRR-!���r��UY����hg�lB(��g�Z�i�'!##����G�e��(j�L�:NL%�b��!��)9��d, "�
�x�/���tk#e�/��6�~<rn��ͦ��*r�C3F�toB-��t�����lٮ��b�v�`�0��3�;w�"�a�� ���-s/s�@.br�`��e2$��%��M���w��{��c�m�@f.�j^����V4An�r��/˳��04�B>6�U���sH��[[�sG6M�W�6�"d��e���,]���<D�^9y�*ʼ��Y$Ȉڌ��L
���v�!�Jċ�l���=&y0�1���~BQ�FӢ�Y�Ya�IÙ��Y�q�<�|B�����D�a�b1uRO��ći�v���E1E�%��F�qHC`#���Ut�0�G�޼�<���}{�7I���ږ] ��s��2���|�Zę�it��a�`B�]�1}q��!r�S��Xĩ)�by1!����I�+���m�~�i/����e�a��c�N���|��Y��8�~6-�hH���	�,�<&��"�ɝQI��dv�'Y�\����!;ZI/�C�G�LzV��}Op���&��MB�"��\��.&T��'$q`�}�:q�!\�����D�Q����-//':�iK&qC�"%8e䠃�������Ð,o�ЅȜN�����j��2�;�S&����T}��H�;��68�(�.2ETV��C��c,
���9`h� ��:@BIO���f�>)M�B�`CDNB����@B�#E*@U�|"'ư���۩��6�S�"���)�qY���������G��ޖoB���Y���QE~�3)���fB� VOZ����}����c�sAXO��K&N�ͅ
3m]D���y��$ G��.B�9�h�p7�#���YYpH���!N\��� �M����`Y����C�bfi�MD���;��*�	�ō�cܔ��U�³0���n$�rX����_ᩅ�20X��W��6�@�u�Wl6�BGrĖ��;Q����ZHo�$�Ț��H�;`�!��H��#ƿ]�$��|��1~]U,=�,K[�e�k���s�����}>/�:J����zq~x�����g�J(/����5�����#qB�!@��j�m.���D�2R��X�)<�FY�ᦆ��{^�r[2>E�H]"�
Ф$F䑅��s���
���1�\�+ɾ�?2�a�+��L��L��t�����M�c��S9R�Ŭ�3i2:Dh��/"����3�L�JI�121�`�������	�
&RR�`������A���H�㦀w>�hh$s���+K{$�=)�*�*�b�
��R9�"�;h*l����LsbT7myö��G����'J2���'�
iXh�.Ҽ����� &�����H�    IEND�B`�PK   sRWZ/�iz$  �$  /   images/750a72b5-fab7-4eeb-bf09-b1fa16e3eb7f.png�Y�S��>8ܵx9�
o��ŭ?�݋�N��(��Ŋ�{qw-�?��L�ٝ�l6���$JME�  �*�Kk���=�u�p�U~�0��u� �ħ�u$�ݪ�W%���gwM'Kw/W��������������U։% �H� -��}���J23�oW-1����|e�D��6�d�$Q6p�|+az���m�';���nDс6���.ǳ	�2��Щ�H �H�3��f�|֜2�.�"��|"(���1�{�r�p���6.����Vp?ᦹޤ'\BAA!�4 ;��q�mhh(��� Z^Q�Z��!hW����㥧D�y+���g��29��8h�mL4D�f��z�p6�c�z��p�����=�h�F!X�T�~�YB�ԯ��\���{|�}�v�]�I��y.�_�p\�Ǜ�b:������ù1ا�����{��O�f�pwP����r�e�M<�������s�gX��Y���D��[�E��;߬���f�qW�`���=x���W�SU�|�Ӛ7��NmןƿK��VOX��^M��6UM�F�(���4��_��}|u�!��˾!�w'��Ȫ���n3&�w�(��K��Vv/c�*������C�s�n���f�u�֚=�n�����z}H���;�<���Y)þps�*��F����������W���z`�9N�=�����?\5�_�M��ᐃo��'f��ft� `���z}�a��4��ۺ���������Y� ���[cA��Țp|Z1��V�J��9��	P�u�8���*P����儲���$�' �{�i�]��1뻛3򭘱)��yM�^�n�ɞmDЮ����o�̀1�������jT�T����{�H�\���׃/���~T݃�k��r�{����=ƣL��H�Gn���ßq{�z���D Pë]ԩb��ǣ�`�v'A�kH��e�l��x]���'��I��Y��;���V��Jxs���[n�F�T� ��#$H�{�М���_�\r �j4��u��u�'Vs������v���ЖF��zΘ۠4���0��j�OnM���k��nm�� ������ˇe%�=
H~�:`�Զ�:BBK[��c�^�ւ�nؕ7�QA�`w�͑	�#�c�P���Z&!��~~~0��p�"�G��k��g������OQ9�N�y��}eDI'1G4,$��ܠ��ץ�����q��xW�%
"��➵ֻK
�/��x:�毵(Q�I�P�K�jyI�b���۠q|�a��?K�����%����;���b��O�s���N:����*��]�2>
�(�n�Y[����=����2p����$3t� ����U*o�Mn�� %f����~����R�u�����B�g�l�g��N�S�Y���ג<�
�GH�w���s����i��W<��^86��/�5�3\�1�Ժ��z��4��,Ӊn�6��DUx*t=������j���>����o�&v���U��/9��q
X���R�"�@^��O�b/��;b����rym4쫥���]䔬�=�1��Ɵ�.�H���¡]��`���w)'5~E�7��	,2#�ǥ���<�@��%p�(w�\�{���-�%�h�~�l�;9�h��� ����V���Z���x?����q�~/A-�L�>��OR]5���_)jm4�]�ۺ'���෮MI���T�o:�7c��!�ʀ���S�V�K���7��ry�=���<Ǽ�27�-(��������Ӝ����L^beӶ��{��Ũa(L#�Y{�GFs �vE ���Lъ������7�vA
�I����mذ�� �̓��|�`2�&e�B���*�V�!������oˍX�$��~�h��-2CG5+_�~q򅘷e��"I<L5�����)%�)�s$(�%�t��w�����J}�p�Gc�D`<y�co��v���h��k,G��y~QTω�`>ԟ��,��3�=�Śȅl����@3�!�=��Y?�'��K/�*~�.�;g�����k��7�c=����$��	 1]re9�q��q�_�MY��] ����Ȑi1��AT:0�_����}�����4�<DZ��r�AC�)�Wu�@��SI�^�\3E�"w!��x����J3�k����a���d�r���3jdL�lԿ�m�Y�:�a�<�i�f�4EE�DF����� �%�����QƜP���'N�5v%�Q�66A'��|)�)�-H���o�8�{�a�6�)h�������$��DfI��8$�g��{�e@ܬ���H�;c0<a��`~ի�f�^!�U�~%�>3�ߧ ں��N�	,r;\4Q��I�Y�W"�9H(�n�w��ka��l	��>����A1� T�� �QB#C�^���8���
����������i�Ꞛ^1&�t�;��
�ُ�iLK��;d��>� 6Q�C�y�Q�V���7�`����BXwW�қ$Q�}���Jۨ`��(8��p%Y����Q Qi��	���/��ڃj%H��2�M��<a�] �T�N��S0a�g�5�=E#؀�I'�r;�T\���\� �0���&�c�8:��Z�l��� �+�&?K��Rt3�/�|I��Fe��+*�����R-���Z)@Z�O	��4��m�S��Y�r<�\�B��fϲ��iF����; ֻ��v��G�B�q��3DK$�윉r��P��pI�m��,�������+�t1R�=���$p�-�Rm�#�B9 !�G2b$���>����Ciz�d2����$R �Qvaef�`���E���8g�	ˑ���;��=�p5�:6�������r��"�Ԍ��԰�$p�� Sz�5���(V����?�`�ƺ�ݱ�R�%�H�X ��@vM��Nfۏ�gX�X��I�l5��.Q�w��ㆵ��p OI���_x���o����Cx7������7e��{?�h����o���k����#�������w~��@��������4Fa��)t1���n8~"�4�#�uF���<(d��)��F����K�;<Qe�n)��$�X�
TD/���K���`���g���P��'04]	p�"ò�-Ob�6��+O���{���}�:r�K�6�p�e�� n`�鯍LPn�I*kRrx����ėe���<�Ĕ�P5L�q~AW�_�͉G�ߝ_a/Z�`с 2E�^�L6��HzDx��ľ/�\\�|���B{#	�!��G�/6)Qh¼����� 'A�.���ԧW�f&�;�E$�k�&|�;7s穽��Z���ވ�o��<ңc��v��M�L�i�T+�x4*Р� �:	0Iа�j`�R��Dʞ�	�
�/�z�^4��544�9F�uw�M�yd��
��^+�J���wg��]4\�`�ڤVR��D����PC�5�6��!'��ܯ�͂�����9�� ��*/���G�+�V����T-.H�Z��D!_�Ԥz�,�D��`9�����s��Hۨ��z��;]���ǟ�"�q���B�W�9��>A�NF+�j�/4�g��΍n;Ø��5GcB����;X.Te�D�ºc��[�S(���t*�~`S�:��D�<|��k���R�u� �����"#u�3]l:�J)؁\��x�<�<�ցq��3&�(���9T��+��xH�#F��u�
��U�CVɀ7�ش��}���H>V�k�1yL���o!J��	)'�ڹ��]f@�˹K�7+�$�a�{d���G��5F��NE��֑dA��5ߓ��!� �؍�i��r7R�˖J�:�\9��^
��T���~1�,�Ј���ٶC�~D��*Ƨ�������zs���Pk	�PG��G��냭MLRx)B�H�ZR�(�ӏ�:�D���YmI�eW:N�� 0y
��׊���6%�r�b�g5��o9�+��W��&f+I�l��2V�c0����q��ڒ��5q�ʏ��<�D��]��Tqx�14u�"B�z!���C��W�ؑ~��熹wj�|��O�AS�ЊC��2K�g����)Pt� 3s�?��@$��aRg�Τ�U"8P��+#�|]��o������t~�?w��vRy�*1��1�B�(��5Fy�D�Mn$I�}y��&.ϫ�3�%���Y��=������߰׫���41%�JS�z�+d���[�[&qc��ϧ����3vUC��O�$���W���
c��5pܢ2N��~�kl凓8y,67I@c��:V��hV)dH�,@[R,����Q�p��߆6��xo`TDU�2#����,f��D_C(��^�铅�� ���7bB�Iv:�Ͳ�_��.`^��|���s@r>yG��:\؆ ��j+�.����TۢN]*֥caQϵf|�.�f�\OQ�^:�IVZ���l����EY-��&�$��	�>ʨ�wK3}h��Y�;�z�4�(x*�D���rf	��?���nmۈ��3J�	�H 
D��ص2L��G����=��D�a��'���:���B�I��>�[�n�K��p3"u��Ͳ>�{a��H�
�ƚ�{oͰ�i���s�Z�9nfX;vN�Iۊ�������s6��d�����Ԗ;#ou��P�{��7n�ݪNѽJ��|���i�M��7�}�Q���>�+��m�9��,�Uɟ�69Yq]{��ryIO�^���_ȧ�7׮.�'��pob�1=H�<lF� ��Ȥ<�v1Z��_�}�^k�B�~�N�u/R�E����9��`&�~��\������u�z�����on:��L��T��G��~H`��u3C��$"]A84#^)Ջ��Ǽ~�<j� ���7��k5��b�L���w��5t�h��^Y�C���'�X-* ���U�k�Qd��">�.ռ:^�q�c)�*��G�P�1WD,ZN?~���#��4���������íۀ�fd��X�\�?��Bn�<k�>d��R���U�(��R��0�h4�"1؆p�ч��� gg+F�ye��9�7��#|�!�}:+?���$~ߟDu�����`���ijlϊ�)8�B�6�I�2,�m33Ց�yn�3�M�d�$�<�(��B��m)��˚���mx�<}�-�֒�������P�U���E?�b��PA�sN\/�yb�!,,�+����3&X?��s�Y�L~'F�|t��^�c'aP\���u];��*JX���n+_�J�谂��ɞ ��y����2O��yLfD���b��#��چߵ�rS��o,�ߋ2g3���� �w	�,#���.��nٲ��	������[&κ[:=���r�G`� �b�x�0B=d��!
ǵ,t�p��J�m��!|̆��h��N�]$M�֠rģ�T�.����Ӡʀ�H�Ǹ�5^�d���Ňm\�O%V�ͮ-:`��B�Xy	v����!��脏�>��"Ǣ��q�vLy9U."��}"���Ez~"���2ԽX��c^�^9&{�hs�V~�f���Dw�`AJ!lVD��Mx	�V��x�VX�/� ��ہ����m��;L�}r���r*5mE�_��B��ق�����
�&�z��Szt��u#L5/L�T==�1�:�>���Ȼj���A ���-�TH��k����䕒i@b�|UÚb[��Cʨw�_^r8IS]?Ԏ��	m�_E�z�=��X%׮p���>�yK������<v�����]Ѷ�G+��0_6�fi��v�DLg�m �����6�/i�χ��d��q$T����vg�g�������%�gn�6�s�_ː-fjw1"���W�ڐ�2�[N��5Fx2�dwb`�4���C46k�[�	����yk��`���5K�����~$3� 9H t���R�)Mt@Dy�G����N^�º�C�y�h���|�j�+��i[e$�,څ���(-U��ZL�c�K;m�2��t"�V-�)�.��SX��
e����HÛ䁄��)�䙱^�!�4/�T;�)hL�.�ܫͽQ��;��e��F<z!23t>���y/�:
qj���8�t{�ej��_�Vh�\ud���J'F�0�R~*�۷䐊��`�TD�Ve�%�s��ԣ�Ј�lvʅ������>��U٠�BlD9���L.��ڋ��N��^�@����c�MO�0yM��Z�˄�S�pև1C*����b`'��=+��}lc�|dr���I&��ekX�7>��_�|'�c��j� ��o';����K5KF�[u}����+�^��d$dd�C?gx5�R��O��� ��P��������$��W]Q,���21����R�=Ռ9,����Ed�����=�r�/�T����=��=�|�[�rX���x�P������a܇U�D:)Y�bQc+=���C�|�aҿ$���C�Y�WZ�J~XE����m�P����lm�>[_�j�r>��!�gɭ�}xO���˵)��6*�p�v���������תO��ьї!��e��$<��y`�PN��Q�7N]I���)��:c��_k?�F1�'<*���,���o�㱤D'�OC��d��}�2�&�As'�s�	�ED�؀!�,~���|�Y�i�w�eiX��>n��?o��׼<>H#��.`+����`Twk]�<)�v�:��{�|u��݃!�l��f�x�)/5x��'d����D�\e��&W��2ً�����E���#�����#ҵ:��|��_���;Yڕ�U���۹J��&7+�b}�:6Ad	6b���`��hNK=�)���H��D��W��鿙M��<���H��$!_��yB�;�s�����Q�v �A����ȹ�X�z�Q��������;䰪C|�)H��{t�@��;�\��V��*h��R!� >A�U'�r��Xon13d�s�޷b�`� E��L7_PZ�M1܄HMu"8�J����RJ�LY�
��i�yf�����9��9c���ҳ��gG������߇�P����π�� ��ߺ�9˻z�C�>h����H�����e�9�}�s�^���L�,�z��a(�;�`D@#m�D&�m)Z�$j��i��vbB��z�R�w׷�,/˦��`�&�i��"3�#x�"J�IW���56��u� �qp��k�S�.����)�vS��"�moe}� ���bG?mtd�-�~N���x6��j��',��f� �V�)�?��W)`{��ͣ�}�
R����DK��R���ڷ��0b�N�"em�#��������79���v��{���,��L-+��S�62�Ww�[�� /�c�����K-9�RUki&��opBR�'�a�o���Bη�i��\�|IG�F��DN[/��x�&Q^��`��������H���$e����d�_$�p���<�`�@�� J]\�c������N�7��	�����E"Ɉ1�
G���>Y�IV�ڷ�)e0*\����Yl5����=g��h��/�cRM�=%�Fh 9�eL�R�*u<�[JM&��T�i��<����
C�ml<����V�R�T�sDD�5kv���6��<&�w	���|�<�2ԇy�j����|t���P����_8���7��'�S��C���q|(_�/�:��Y�n��ׅ�[Ь� ��F'�ĉ��#!"K҉{�63͚�K>�����VD�2�Lq�S�����Y��r���?Ϯk�5��$-od@4cvP6�	��ܝmX���L[l�o�/K�-%���K���HK�*��ny��ޚ��n]�n����]Hib�;T����s'�<1���{�L�ҵˮ1v�h�C�g�Z�INُ��D��������>��w��E��'
�<]���4�a$�SP�q�
;TE�Q4f�é3lD������I� qü�~��g�57<�|��жt�4�d?��=��8G���W7~��%[y�g!r�*�g�:1��7&��}�+�j������	���f&�weO
�jYX�U���Lӝ��騂��^��I�V�.��P�p��0Jِ X�K名���@3�˲H��Q�R��Ǚ�XGT+���i�;��?��)�[�"��#~\q|0ϦY_l)�k���wN�B��?�;wqM��$����ƵNk-������������He�
���PA�P��h��a�2�,K[
�c)�k}�tɫ]������.�B"[��mp(<)|��������`���*���ӄmE2�V�U�K�� mL
7L���^��fԉp
���y�iP��+��j���H�r$HG�qq�Yq�~bbE�stM������ȟ�O�ػU�T�B���фK,(��%����d}�u�����aO]�N"TlԔǙQ��� ���)�<H�.�/%z0,�1��Z�ҭk�c��{1_0�.}�?��T��wzVW��EB $i����~����q= ��\�S�ݹ�2�j��l�K�B��g�mX�ۋj�(�-���F�>'�s��W~eg~�.)�����-�mQ��I�+�m�b���=�]nV��v*��S��9�ߕ��X���|�(�8��:��٣�����=�&��ꄜ�����$[*��&�[i3��bm��t���fxY�r%#���`�\�p�"a[4���D9�M?�T�^�������ݚ��,�b��p�(\�t�rf��+2��r�^��d�-Zw/���c<��u��/��I�h;�>�!���P�[�I�(���Z�B���ljj��h���7F�+)�#��%V��:���]�E^3�?�8�Ao|,&5Mm�Y	
���Ͼ�\\�3!j:>��2��S�$�&��m��6y�?�s�sJg2�m�v�\�����O=�I��������]4�U[�3�V��&�T���m���VA"1��[ </0=l��c���WD�Y�٥ '��X�s�)w�D��+9�
�Ж�֐f�|M�c�G�RLKy�wWM�H�3��Ϫ�Z��A� T�k	�P��T8��HN�oS��`�zNIc�<��6+ϛ��;�����k���d�(��Z��%lllBΦ��d�g{�8�*�s
ڝ�sg����.?U�iO��P\)�ܕ9��Й�T+��1{%��"��@z���dT�+%���PK   sRWZ�Ba�  �  /   images/8da9f3e5-57f2-4cd5-bbab-5c1279684e76.png -@ҿ�PNG

   IHDR   �   �   
 C   	pHYs  .#  .#x�?v   tEXtComment Created with GIMPW�  ��IDATx��	�e�Y�y�}Kf�ܳ�*�-���RI�eY���0�h�=@��v;A��#�a z`�,��D�FL0�qm��ॽi��*�RU�T{U֒���{��}�|���r�LUi���H��|����o_�_1MSwu]]��J��F�i�h};��GQ�_]���؅/�����~�w�ԩ��������G��K�z���e���/����"+���Q�1�ԥ�}�ꍆK�K]��P(N�����P�]�k)��d��κ���Ǧgf޸����.��.�#�rss�������^�s�RiUWz�a�����w���Wa���3��$5-��b�認�����Ca��&�&��Ԕ�׹�9W�Ք9��Z���s�S���s�=�n����^ggת��*�\]����IDK$I��T�8L�$5e����'''q�S��(�nbb�]�xQ_��W-��������p\��Ԭk��*���7�|�k���8v�uM�2��u��c�U��Ƙ�I��O�V�w3�z�°�fa�z��yԌ�AxM������j� ��X�$��0ׂs�=����Ǣ��q�?�*ül���+�����P��[�Z�.(DY��/$"�kB�����9��;	�ƅ�����]��.�N<�N�8��Rh^!|��k�H���Pu����J��9�&���6�ǉ��z1���淸{�/�����ڍiڝ��u�a��K����6��T(y�"M�� �B���"w�ԩtddD5�����G�q��������?��^p��?vL��w�OU�M#�gE��w���ÿy���J���lbjl�2JA|c�n�A5��^���[N\b]e��+�6��FRs��`ɓMma3(���t�sU5�Ν?����4�Y ���!�~�:�/L�C��>��j#�ʴ��t����0J&��ZI��8���|�o�aJ�����u��z�7���neԞ��i�&���놆�E]���=��ܺ�0���L��o5�tnn�cB��
�+�l� ���1�3f]Q4II�kJ��7|�ٙ�<��[�v@��9�����3h������֦�]�|ƪtw�m۶)S^s�5��[ww����5T#6�����i�(kۿ��]��0s>�̖�XP��h�K�H(N��_�^�nm��/D����Ͽ�����|�!_�L�Ǎ=�B�j	_tv"ջD�̹��Y�n��Z�h�z�N��L� 0��[��߇6lؠ��V�h�A��nܰy�0�~�I�9E:��6,�>p��#V͹�>J����a�,a�b��*L@��m��8��&��ZE�\Igf�E;��8+&Ԝ��Ը��)!�9h��hf��a��D��p�1�3���`0L-h�n!~�Sx&AS�w��Q�7ov�ׯGC�!�0	�O�Tz\^���ۻ�'h�����D�1�
�h��̺T�kq啌�53�i09�	�������錼���bͪ��=#~��iӺF���X	b��,�F�����["!H͕�hvf^�Y�5�e����	�%̀���L!�﮿�ze����s�4�1�|�>����{B�A��w *�t4�RѮ���2�Y�,���\��Z�.����a���y�������6�C�b��(C>�(�xa�s�GU+���l�ʈh^�3�7���ɚ�̰e�V748�D�'L+~��E8�.�%(��:�Q\�}#�����s��H<VUSq�0���i�W~]e��.��6Fh�|#q5!�Ύ�p����dfQ�E�\E=�f���5Lm?ih����nttLM(M�}��qeL�7#��JF��Da���&�5�F������*��p^����7<c�\���̰c�N�30�zzzDcL,k)c��l�*�S��0B�%��w�m��3����[�7h����`�U�Ya����V"SM�/��= �\*�����SW*��K}�M�R��߮{� ���1����<yB�ڂWoO��z*�GC��|��r,L��������
s�%N��'	=q�RG��&�x�!|XvP��۸i[d��,���.i2la�������*Ä���WQ��ue�{���JsZ'	Q���B��dO��:�k�R^'�'�����*p�D@����o�%��^�ޤ@6�Fc�DS`��=���|���� l�H�'�n����h�k��VM���'l��h��H,LR�����֌y�3�
��+��=�0�� 3V����=�q�'��Γ(<�B��I!��A�����OL�	C��[�������Hj4F=�\g�Tvqo�� �{���bB�9e�@�%�j|��k0[|�i�fmq��s�|����R��1]�����L0%~�(j^�5�}������z0�r��K���B�4�M�5�_�8><i����H�ڛ��44�v[GO�~�ւ8���Φ"��H�ibb�c�Z�"Q���D,�Cפzwg���Rr~�S��ۛe3�ԣ�����a�c	@�._�(Www���+�?QQ�زy��.f侎����\.�q�0i�ig84����y���cmH�?�̃��������n�sl�}E�k�a^��u�%D����1	6�T�B�O�6~�f�e���7LM���腇�@a&�v0����?|��x��t���sc�c�ĩ3ZB�)��:�*5ܙ�g]?�o���|2f���kU�����C�96oަ&����ɂG�v��^��������e�LsED�J�X8�5u�+���?5>���s3�W`>�;;��{ç��H�2Z����%�]]n!h���	W;r�M�x?q�8�]ndl�U�*��԰h'�]B����4F��*��,"U^s�T{�tE��H����jTj׮��I��D]ݽ��PmѮ�M���\�g���-V�������zM1̕��J�R];3Su�c���������;��aWM�0?-�dF�?�!<"?q�*"勥��m��p�e��0�Μ?�.��*n$-���YwntT�f�	!�����qWr�^�+a�`R%.�r,��`�߁�Ŏ;�u׮��o%�!>F�����-6r���U����c3�g纪E��z��f%Q��yj��� �-:�Đ����M�T��#�S��p�a�ӧ��ﳮ����,�5��%NkG1r�R�:*.�N��ܤ���R���*ٹ_�T�z�svv�97���\��!ڪ���ܜrT�묺80?<��/��j�n_�i�F�($lKtJL��{{{�<��z̵����6עHV;�D�K���􇖲+����^���Lƾ��\���0>���`�Ց�1��NyuN�F��z�>|��"�
shYF�*<UwgŴ¬���qe!P��sZ$�s�5�ı#n�6��&�Y�����P�viM�M����D$R|c���:+]bb���\��	U1��\#�d�\�r�w��������շ�3����o�~�0���1���wu�6�k�a4���Qlx*f;J�	z-FGG�g�BI9��/�h"��=uf�5���3M�6A�/�7BmTꊱ0AC��6�Ra�H~
�+�U��)�MTs�hA!�R-���P5W$X\p�׹�I�+u	t��-׺�7\�6o��ݸ�u�;����z�3k�J42�"����K��o�E������Z��z�&�@�h���h
Sz�ye�b�}��+�1}H�4D�(5'��О�j��'Nd��Kcu�!Rr
��gAL�d^|����y6s��˩�)G�8�99v!t ��V���(i-��7ub��t����~�K��kj��}���_>�JqY5�Jeb3#�	/��j����1LC��"�5���j����N�r�YJ�Na_B��!�E�d �S�Xk�Ify��@vթ��L��@i�j�S�����[�s��nq����-�n��)�A�mW���$��.�H���(Z-.w�s��\wߠ{��n�]���kot�B"�K�#'�) .6 ��/#�C�R"V���%|�K}�_��X�z�F��?�Y�?� ��G�U_�k�H�I�V�B��W �����5�t���kI�=���P
�/&\�U��;Kuw͆M���¹��̎�����SpC�}��j��|V���(�$�+����1��G���W?����pO;D
�Jpߛ�gsla�ő��~�i��/}	���4�;�a�&
mAC曵��:;������ӇR�n�-&�h�2ߋݽ��톆z��-+��|��� ��וv�������H\�C̻�Kع�cR-�F����� f��I��#���c���6R��(M[)�$�*�,�B~O����U3̢b����Y���B�ݢ>{VQC@ټe�f��Ѩ�v�3���ū-$>NyF",�a�&y��֯���޶7�a::J!�
 �0i$�J�D�nbB�~1�:+¤�7��h���	7=;�:;��+�m6r0<,"w\�Lu���s��7�|����=�f�m�-�}���cw+{Y�׹�����Z�(���3�ږ�,���R���.8�e�7|��t��۰n��3)�7�������n��Ӝ���kc�к�O̭���X�1����"y?"
=�;\#�G|(�i��[�C�`�ti�H��=�2��N5��4q�E���+]�v��x]�7���E�1�����?��/�nW��k�>̺}���9q&��as�F�Z�MP����e-��
������4�i�vI��Z���ɓ'Sz�u_�u�bVAX����~���T��a�	�b�3���'n��*xuR�s�E���;iQ3��ǹT�^�\�h1�f�&4"7W%" �V-tOF��y�ɔrh�q���-��7oqE�^΁V��L�`U*=bnN���>=����m���~�~�V�[hM
�Kݾ�׫���3:z1>�fVJF0� [�������ܼj�RG;Pt�Z� �/ ��l�����oh*=�{m������F|ҍNκ��y��iF���t�-�43��i�*��H����U_i'*�D���������߹�1؊��m}��w4`���6��E��Uk��ʮ���<�����|�|�W-J���|U� �`�t�i6oޤ5U_��W�}w�������H���z �@ӌ����c��@��(���А�P��"��/�����]!!?����UrS�5'֟#H�h�{A^��_H�um�R-�����Z����𘛜�Q@���9՜�iϸ��!<������மﺥ�Q��f�����>�?v\3��ŋ�-�pWZ/z^�;55��M�U�}}=ntlT�	�!��O��Y�7Пy���"��y-jf@o�w��&�E�ܽC�d�IK�c5��3u����u��dME��t��PfHɛ����k	[�Ţ{:N�W*������'m�)��7�{���������������b��̵��I�^�����4=#�z+Ŋ:��W������{�ȋ�������ٹ�`�4C�IhbJW��"�W��=�pX��T�K�h	K^�W9s�LJ��� .��h��CTL"
�����q�5])-���j��$�e�{�j&	͂��l�Bf����
��@��_��۹sg���F0�^(\��7��a N�����ϧ��k��N8�$<���A%f~�J�!�V�V�I�>&z��U�6����caa����jծ��1� �b�Y���.��4ñhu����B �akL����4�!DF�OR�lCh?$+[W$n�̢L��e����h	�\��TuQ�YO�<�Uc�)�����q��=��s�4{�E#����a�\����&1�ȋ���I��"�O�o�2ؠ��llݼ1D�|����3�_bb�����{�{�������=�֟QZ�R?0��;�0Z�Ul�4�9�>�ң菢a?�^�%�X��r9��3H�T��z��(��KH�@�hџ���w�w��ڵ+��a�;V�0�Y�����C��H���p��D~��f9���͵�Ʃ����KW�Í���뮻N;q�Ak��U�uH��h�������=�Ѧr�GFL2��<�n�����W���ژcO�т�=%M���j�M�6x��0sq��h}�YnWX��EK���~������V)h/w�ޯ����)0l�[��C/%ڴ'Ey�k�/�Gm�f�r�ɩ�ӷ���m�J��R���2hՉ��Ѩ/�l�a���i�~�y>�F#`O�s���_,���a���h���{.��t9��[n�E�I�+��I���I���P��!�	@�qt�V��t	e���j��Z�]�j5�r��te'|������������AĴP�4K��Y���]"��?c^��D~�����n�~�4��	��A�������D� l����(�ՙ�����.Y���^���x�Ϟͮ3�0ݬ���4�}��}��[o���Jm�}�}(�l����H�я~T	��]t���faf�	�:������L�_��cƠ�ؤz��ˮ��X���rg���襯-���G�m{oO��K2k_�RK�}�zfo��Wz��%BW����Y!�����*"Ε팄��ё�E�e)B?h��a��k^g�fL���L+������g����8G#צ͂N�� �Y��CQL�&/��.���G��AK�g~����-3/A��*���?��zc�1i���rr.�<� 4hS��}4���Ѭ4�Qo��^��� ˠ�WumٲE+�A��w�?����=��S)E��%��:~�x˿G.��_�`�B��aډ����������"z�ʞk�����'�/�wM���� ư��ZJ�����c�&��� +����D���g�2�L�L���IYNd�X� )_���܋/q����?���%"8e�&�7�쀟�ԧ4�MS��_Ka}��Ϳ�7 ���������{���`/����2�*�:���T%��u[��nR�2���}��>>�s�3�|~1lU�V����J��_6�ƥ��+q�+��̙��ӟ���䣏��uC��ՄH�?�/&Q�x�Ko��(�k�e�	��Β�����\�}6�i 
4���	��8r-Fd-�Q^��__|����M��?�� H}���L�(n��u������h��T*�Ú��i��������~�1}�/��7,����	���
w~�2ċ��)T��I�����!}�K�I%������4��x��9������?c^|!A�v5�֕��]��D�̰�7oڤD��a�P��o6��e����i� ��_�{4���R�)W%m�Q��.e�b�b>]�ۯSԹAR�c�F��=��M��)�%�a�@,���/��>�5qQ8��'N<`"5 �|�niF���ꕲ4U�I�øּpr�H��_�z��H�(��\G�iz{�3�����/�Wre�w�Z~'"h e��9�]�Y(-`0�x]�RA��ɳ���,j7X�N�VɟC
�%I}�8�\�"�KdO:��{ќ����71�q��Y�l�w���I9����>�������V�9[E�h�~X���l��=�jrZ�������@��y�)a����u?��vO<�D��&r,c�i!�$Z�$�_�����|&��Q0�XD�0��}�}�����9(]H3�5���*Bɱke��t�����`��t�����F#�KdZ0m�,w
�P��~���}�*@�D#+>2h��h�  ��߿���I����F�/vuv�s�Ω4c����m�'*���Kt_���@�+?���%/e�u��ttt���Y���py%�G����G5d����Q�7�&�D	M+l��Q�E�V��]�j�DK�����Ț����5�!=1�[�C!^t^#�-i�j^�@H�՘��"`��v�I���)魊z�IܦL�{�u��{3�c����(.��Ө��ju?���P�e#<�Zs�A`Gix��^_���<�ɱ�}�Y���.k��(��6өh�l4�юgO=�M�l�Ɇ��ry���R�x%Ŏ��.e��Ն�+��f���v�$/�e_��g��~~~gR�w�9ggZ���`@s�m�F�����,�,̇/|@!J3�^O|iz���Ʋ!�c]/����׼4��(����DGĉVY� ҈@�q�I���d&D����/�<��ԯee�j9�h9[3]	ǘ�j%.w���D�K���%����1�ɰk�C[�3���=�<���3b�L��R!�{�HCCC��4�8zR��\�r.y��O}�,�� ��Z���͉g���������(��i�錠֭[�=-S��;�Y�.]B��K�ſ_>��}Ǯ���}-�/�3����T���~�y�vӐ*���ɿIjC����]�i1�i�h���o�x������WӊJ4��{�'3w�%\{��	a��axs� 
m+� >&������t�$5��k3I���q�S�ER����8�J�+vx�5��.�)�)%�D� �8~꤫��R���{smY���Rk��	����͉^����� ��zMSΏ� �ߤ�H�$l�tܝ�����,w��N-�`�f��+�����OM����0��7�H-�g�� o���-�efs�xY	���Ȧw�u�۵}��ޠ�����,�!����:����GC�T�Sֲi�&�$�u��ϴ��js���������E���8�v�����/���{��	����"�Dq�rK�M���u+�<P��c�0�Μ163��t����u���F(�,��0��z�����.��G���u!+�9n׃63K".-���EӒ\��Z}�������(�8�WB�qaE�����=����>����[d0�ݿU��x^�I�Ua�`} �׉Iu�칖��tXnx�:���*exx�{���]y�#����J�\#��ܫ�A0�H}����3l"T�_��a������,�0+=d�>D�4�(��n�ϡ�����$�+H���Y�Ԑ��J��A�r��zy*=!m��`T���f��43+���^	0��S4������r}�����**pTaf���dp[H�{�:���4��G[�_�Uy�������m6�×�P.E�Q�9��b��c9�����f`��L%,#j����X�s�at��ب>GjӠ�.��f6����H5c��%k~�U~#�3LB.��d�1�H�x��(3��>�+T��i�������@����K"@����ucc�hT�wL@E8vTTc��+�,�"��n�:�m�����>86:������=\!��%-��&@8Hu���p��e����|��*D�L�^	���b���639�&Y�T�W���h? w�Mδ�啞^�칍�RD�0�Td���7�qG��E�(�d�� �hX0��4�t�zue� a�����K�{��7�oN7)�	�\����+���3��:����~�J�ut�6��r
��ssUE�t��)�`Q��Y>cҢ�����*�W���U¨�$��꧂��}�ww�~�}�_tO=��0���pl�K�@7�����zk�u|�J��q�.��w^���W��N�9�ӺW�~�uOs:g�ɹvk�UEp���ՔQ���Yj��@���~�z�ɽ���q��į��JL=b�)̔������0w���g�m���~�����3�a&���"]�:qZ�鹏��v���/��>��MMθI��b�l������S�ǹ�ywĽөψ��*%0Ȥ�����Bm^�=�
ъ�ͨ$�:=���g<;��{��5�r�r-���MY�af�m��N��ok�Y|��K~>��C<6�k׮�IP�c"5G/^�v�|�#���s,�E9е�v�R9~옶+�9�	�G���@�H4*����.���05�U���0 �����v7 �3,��7Ptp�i� ��}��
�[���o	o[�*n�9Wby�ITˑN0_vLG�$*�|�@C	��nC��[Bɻd�1�J:1Zi��:=�Z>"(1��+�G�����z�9f�KYE���ǰ<J\hGb|e�営�_��!�EI~��aw��q� gD��C�|�w�}�0`�DG�`��}/�T���?����P0�A:!���w���	a��'�v�k�f�\{�2*��"��B�\6�1/��k,$�|1�O
cf���Q���\��Cq�M7)�p?|s%�L��L�.�7�|�G ���@��Z�q�w�~J�N�8����)a��F��h��l�cҔ�R��=�nI>K0_��^$����0���	�u-�0�S��f��eK�~�'n��r��Tۙ{@�`#��TTL��\ԁL��C�H.^�C�(��	��F�:4*��f�yEZ�=�= �H�������hy�7m�j�ֺ�`a^L�c�%8'R�J>,����� �lhA��!�R)��T���B�|W�B�%�\����|iu%�]�Q��׉�fq=f~��1���q�d�y䄠Ĝ�I6��!�"�5aLXF"6�*L�0�SF�VG�Kgn@	A��y���p�E~��W�w;r}�{��Yu�2߿L'ӈ��	S��|��ss�S*�݌8��<s `�̟���z*Ff�S��Dnntt�%y�ԓ�R�"�A���5��T0%���Q*1���]�ss^�+Yoa���z�6'�gD@��=łZW� �T���26�x�	�v�A1*���!R"R�&��<�R�߾����<BQ)���乨6�'�"�/U 33Ӫ=���!N�<����d���(��{�tu���Y���g&5� �D���)*$6�Q@i�����������6j ��!�����VZ��HV_����s� �&��>���0}�H�����yq:��$ӊ`!@"L���Z��I�k�.�������Qo�լ����|��SH�?п�`�+3�亐��߾/�_��/?!�T���s���m�I����'i}8U{>J>���	�����1�����Ҧ9��ъ�pN��v��x��ôf��>�g�d�6��f���lРh��ED�:͇�I�������sФ�!���h�ԃ[��[�5�kkY4h$ �0�>�����u�-�ܼH6��iY��|* x��T����N����^{�~�����hŭ<��\�?�_�Q��j~c9��L���[6o�(��'���ϸ�`�Z�ܣ��#�Eu�����%�e7�������A�?�Ϳ���9��
X"�WQNҚ�h5)���\h2�� 0�΁	��a|O��<�yp8����Q��P��AU����ѐ196L��gNgm���r>�b��e�{��&ɂ��9�h7����
M�#d�V�>��h�U���_Bbl�E4�P��%anV��1��	�]�����!�:��H���40����7o�"��u*i��}��^ �D��g���+-�b%(�HN�w��Q �����ֹ]s#��� �0)�Z�O�N�Y�7d��q�������?�C j/�}�Bd0��UZ�ɕ��
w'Z|J�{���'�s�ݰ ���=������-�h�3�ŔC�O���^	^ �u(�U&0Z_O���a������i�0�O�pOOv�V���+�9��48���щq&�&P�Nי���_���yШT|�F��)(a9�,��V����F2��L�z�{�YRm��*	�U"�<zR%��k�+�oڴE�h�:+:PvfZl��Y�{���a��l�r'66�s�#Q $=��Q[�&��o�j��ǎw7�ޣv2��Vç�1a�3��z�R�����ug�� ���ѣjj %��s�W�a��4�]��+��u@Tֆ�y�D����	��!�C�:jk"4�m���+%�PZ.,����x`V#�U�����a�}����*^�oߡ���,�J���������n
��t�0K���	��>����%�H�$`9a��]�]n.�;����j>x��y�Hg��$���Er�^�!�m۶��{RÇՀ+\��6�sAI�eo�CPHn_�Vp��B�;�z�<�4|���`~� � +r�b�]�XP�N$"&e�0��������p$L��̵�
�ɅlݲM$��<T��566������/��wM���O9ج��9g��d�=����+<���|,%am��@Z�i^�k%"o���Y�H�ߋE?��f���5�ǩS(���U�,z.D��qI{�3DQL5�)��|��	u���S%��^*�тj�[-��,�E���R���s�5_���"yȝr6|��nQ��@��n٫jG5{��9�Xfэ�^���S{Z$��K�,aZ�f/�;���W��ݻ5��ժ$��D
hf����5(����Cv�ɴn��f��<�3
	Q;��ވ,iF��4��Sb?�>��y�F��`4
	7B�|���	��D;�o�P���'Ab�/��y Pq^����ő�K[�(���gf�GY��i�N{؜н1�W��ʁ�,#P�%�dK}MŌ(���L�s"�i��$���^(d�'���R�>{K��9�EW�Z&υD�$�f@�.�y�4�:L�>�`��B�"9�jn�eO�$b��r�Hf�T�d�Q�h��E�#��d�1��,2���?l(�Ɓ�9����`����@�t�
��(�����p��yx��e�>F�`�9�'[�wQ�̞8V���'4p�Pv[�nՇO6��G���u����	08/�<� vJ>����T&���%S�4�
�'[�f�!�d^��v��̛d��}ψS�rW��̪�\Ԅe����~y�zJd(���y��ξ"$����e�|M �g�`c/�g<v옛_e^&�R��R,�`�af�;V}d�:�%	�b�}	C�������=J���VT�f�%����\�蓵�w��	�[|��ϋ$G��^�ZA��2�!��ec�/��c�r2<$�J)*f���e:꘸_B�۶lu;�ݞ�������*W�]Ӧ�XM�X#�~�1)�vw���t��:�c��MZ�300�:�:��"FyZ�i��)��+wtbQLNF���+�sZ'&#�ĥ�J�g�c�����d����yV\���XRT��gg�p�]�mb�~K��'��)�C�|5��5o��aN��<IⅢ�*�Ϫ0�NMs����E-l�����4�x�3U����sY��ֲFr����-�9Pӓ]���s�7g����Yз��:���N۹���cj�hFL�a-�\'�����fwJ4G�Z�k$¤��M��l�@M: �~��n`ݠ8�/�Y���w4h�|G��w�¾7��:���d���j�@Z�~H�O"��={�3�|��'N�TP߫�*�Ð����\��z�K�c�)�B,�Z�P��bA�o0=R��>��ZvK�a���/�o��}4�Z�{0O	"�-̫Ƶ*k[q�o*ľ5͎�Ɣ�/(�-g�|i@���~���n��>�^\.:`�w�T�d%z�bCy8Y�!$��[TҪQ��U��w��4��gr86A�-�B�6mT��=�71S2 )q<��ΐ'8191�vl�����1�0��H'�3�:2~� �&�衚_a��Bh��U3�G���T5�0����y���5T*Z�����3�I��!�B(mB:;vT<�	����)	��
!�x~X�� ���`��_�C�W)4yY!��zu��!]�ÿԪ����,��/�4�C���x]��g�����M��f�)�Z*Bf����1L!�YL]	?n��������� z����N�]����`��a�ld^~�-��<�r-�v>?,�#'^j�_���Iu�{{��적B��P�G�Ph~����6�m�Lk���=L&$��7�Ԯ�M�j�,w�y���k�D��s#:g��#\a�J�����0�p;>�@�Jh0*�#�(6?&*��s^8�]�}GV� C:?����7·O�J�ߓ�X8���&�K�TPs]~0
�ڄ=ŗl�(�t�2���:gr�4�_>4�bo���Z���̮�w�̫�������1 �:� qQÚ�";��z�p.�܂5�=?�Đd�o�V����YIBE.Kh�Ķ;�ɿ*z	9���ħݒ�HI}a����6njD/�M\+9a��&��Νvs�t�����^� -c��c�IA�4�腸��GG�K�Ec�R�\?�/��L��l.v�������|����naj�#��1-ޔ�b
�_fJ�[�`V�Ǳ�'���_�#��t>l��J�Xʝz�2��R���y���$�ϗ���2�ڂ� �>&����ɝ��zؤiO�[-�Kڜ�����q"��U��K��(��a�Û�MX!;�����z�hO�U�x��}{ou�Ť����Z�VHk���uWZ�HkV� �}�H�B��ԣ�42�5b &1mVK��-�TrC?����:���"��7`�x��dV���D3@x���VŢ��C�H�ި/��0��R���-A�{ag���Ն:�����
0P98��rjݶ���o�"�j3�Z9���;�T3G�1u��~@�Lf�T�t]ͳ���Go\j�="��h�Ml�cvv��Y��Y QPɢ��VK��lF3'�>���f��"TK�%l��H�< D�/	!ClMr �	�m��Ֆ�7���4�R�&aћ&����%��u��l�e6JaJ`�sB&�a�7��
�i��F��E�b�@��U�<گ�����?Z����o��e)�w�s �5E-q���Ą����&>AA��,�mu^�������}��P*W��+���e���/C�f��P��Y�0t��4?۹,��~}-&�d j9����L��;���	iF��8咏��xHD艠�qg�-��ܦ�f�R�<1�R-�nggA�������z|��zF�x��I0�5hL2LL2�s��-��<���A��B�u�8��18��V�(IO�x��j���Լ3[��d�]J@���Rg>�h�Q!G�oIH||�Տ")f�Ӵ���}�j�	��+�d�_V�R��s��/M�V
N��v�'c��=���&H`(��o�����BM�y~)�[0�}vz�G&"����T�Ckj��..�����K��Ȓ^�<�շҩ���o~�JZz}������So˦n�u¸�u$:�r�bv�٣D�ēO*����ٯZ"�(� GuǾ}껠5U�ʹo߻O���sz	�o���ࡃ����M�7�׿��Z^C����{�q7��E-(\hi	�StlzԽ���4�A����N�xĭ�}��-ʔ/�x㍊7�s��$�I���ve}Br��r͛4
ȳ!��sܿ�@f�ܰk�V6O�R4��s�k�U[�n��Z�{�{U���}�+�K�w�j�����p���RQ�$��J�V� x	�N��	ݱ���ONk��G1^ޚ��R��9	4h27iPϘ�z�D$m�X�'��ʍ�Gɐ$ڠ4;�&�}�n����~����L,��n�0�4i+�YI�3m�W_LCy�5̈́,���!��)��<�?��!ޱc���@0T��q[�lu{��䮻�,"�/���T��0Ԙ�T�|ꛊߵS�uH��ufE�jJ�>���w�����|��l35g]:fX#87�I�O<����觟'��wܡĊ?A��-o~��B(a��z���zJ���4�^ ^����������G�����U�"��a�JJ��;�|�o'�������7oޢ�p��ݏR8�Va\����B�*�{����@}J�ך�c�����|��H-��4]��7�~n�e��q`�h��8�����i ��
����_->L!��[j(���p$��g}b�%��ۈ�q�]]}Z���9BD�0ú!�=�ͪFڲ��C�)�B��S+d�Kj��Rnq�o@q$e(Y�2d�!�O|�� 7j�	Q0��ҁ���b��s�Ѽ��q��Z�p��� h7�}P�^�>�� E��V�n�
��=��� ���I�y�%�^��+��&� �� #@ܿP���c?�cZ��!��	w�h��~���_o�;܅���?���=��Y�{e6
��s��|K�hȓ�д�04��]�(H�b��8�h�4�b��F�����>	g�����e�Z9>�M�؏j�3��JW7���ۮݞa�)��U��q\pǏ���R���4��Ԣa�g)��E_E�F��&����^���j�hd��:��CY)5�e�&Y����xUMw`�����B$��l�Ƿ��F[H��l�x��b��v�R��W��Ϟ9���[�߇Eh��{k6�aj/=��y��ӎ{��ǲ.������36�^��h�{��/}IM�<@�:�i�@�hT4�QU��(1r|B����̵�|0�%$�y�$)�c߾�B�ڗϳ7�H�ٵa�� �w�}��_T��7�I��(j�S��z�.�4��9A'�Q</�"Č��b�;׆��}�c���Z֏��aR�1��QO�G����~�t�s&�\#uP��"uD�0�Y�bU�G=%����t沟���F��]�0��|A�V3���\TĎ��(�I���{n�lYr�ZD	�����3"�/�g \�l5�t��K � c�G�嘨}��i!f�v��w��>��ϫt�����駟��\��k��j�7���A0�E����׫�"T�a-�B(���>&>�q�D�6������#?��*�)-�<�����\W@CyF����`k�^���o��7���c��gݺnx���.4�����5����m�����,�j]q�DQ�;ڭ#t�z[ƽ��oU�v�MYn�^�5_��Ν�<rK�:��)�ӠA��~ �D`�@���N�l�(צ4S�=%wͶ��ubҡY�.s��y�-w�f��·�>��*�RWY�v.t���t�R�	��;���1�����������i�LlJ��0�V��A�r���7�}�2҂�s�i-�i��lk�ȥתvy������sh�/T�a5����vHQ��^�g�=}����Hם�v�ĭ
$*��:1_�h�c���	�fm��y��)�LH�hb�lr�J�ݡ���"��d��͆;�� 6?&#�6_4Aڨ0=DcQ��`����>/��^eb���WLK}T�i-3�f���.%o�a�l�L�z��Y�7�� ��%Zڄg����p�[6ou;v�T�-�s�3sb���]8`r�^(�P�m����������-ά|��q1���n�ejaҐ��>�'N�LL�h��{��Z��𻰕��|��|[j�7H�u��eؽjr�P녶��ŉ4�+`8�H�d�ђ��2��B:�������%���Č�s�݋o<�}p0*8X`-���i�+�q��S�%"Gg��m�6վ�����]�5'U[�}'z�o�F�D����3;�k
��n^	�ɗ�̫6ޱ��!!����P@E�aH�
��}��(t�5�U��UD���hYo(���r���Cm���a�-[6�s߮�J�=�� �� ���������`J�-I��؄=�9�2 ��6��x��w� >Ѯ]Z2�I�o�͜��g&�V��S�! ^`W��ruާ�|���*���]�A/�|f����CR����)��t������JAlS�
���svߴ[���3j"h-�(����[����I8�9!L��S�!�q��k���`��j���0��\cs�@Q�P#�bfp���7�B���(�z+~-05ϓ(#~��ۦ�$0F�10DC��,��Pԗ��0
UA�m��F�E-���i0�M��ܸ����ӱ�!�Toc��U�е����q���C�y_9�c	�}�qp/xV�h)���\XE�mr��X���V�0r#�v�,<3,?���ʪ}���'VpiQ����B�n������&u�F�E�F�ظ�E���ח�����Ci7�y��K����7f�{
~����f�sY�	��}�ڵ���&�&��b?�8zܝ[�0�?�=��l��ʅ�#Ӌ�� ����� &�U����Gчn�&0��oݺY��٣)m�(��>p���H����g��LκI�,[6���ة�N�� �����]��'������@J��a2�ɡ��	xd�� 1�?�g=�H<'��z��e�VXD�s>?u��`(��s�9���7�}r.�"��B�bB���� �㠁��F�ߍ}���ɓ��}��ϩV�7[�q�����.��gO=��\�iը<cLi��4�4�z�Fc�d��}��n6��_r!�9�lHs�HH	gΠ�L�O��5_�w�A�G�U�g��Hl�;�%�$�6X<�b���T����>�Kd�(
��B���׍�j�U`Zq�ͦ��T�����u�!�*���0�ʫ���P)��y��r��Q<�2�`L+�۷W��d� ș$�ٶM%:�*`L�D�t&���Q�&g������'!���N&�\+�v�-{�����zm�*>���dD�-��bh�C8Y�F�<ڨ�>'5)����lI�R�iv+�/3߄D:�A�M�z[��޲���T���X=��hYm=A[)�QSH6�j
3��y�zA˜Ȟ�#�*��0��z�������J�Z5 r*%u���2t���ǭ��7�#U�΄���@m��l 	FN]~��CS� �'R���D�a��Y�����,�v���p}�� 	����g�DS���V�`*�Q��d���|�r��MJ��Ay�H���z^"G�0�Fy`�vX
0"���G.i--!*�k<p���D�0�S��7赐���w�@��~Q5���y���{v�l13�`^7mT&�r�b0�B��0'�	������#w��y����h�����:>K%�����>P�D�C@�q" �ѩ֋� �B i����>�3<h�Mi�V?'0t���NJ<�S`
B:}�������낯;B
��~,�h��6<���T:�͡�k�4��z|���{�I�zN�7Mrbc�
l��Т�[
���-�d�����yES<'Ďiy��57��ۙ�a�ǡ�t.�YB)D���

2� f�Ўuuoy�[U��ں՗�pN�Ï㮇��b�5��L����#� ���в9�������Z��@�|�s����'��Z0a!$��^r�`�i��Hx�z%%Hl�J�5hC�A�0\�EB�D�JRDM���46Z�Sނ+���� �x>��{a�?2�C��/Բ�&�h�&7u-��$��{�M
YˉVo,�aX�f��đ-��O�5֯�$�!�����:�Q����wU��&,��HQ!j�ņY�R�C��euF�'q()℉p[4��삖�������Tvu�����U�8*��1��,bF����0�׭��r��m�>�暭J���ӈfVD��i!�a%Z�� �@�v��i}�C�S-���ܳ������C��D���>�p��)�%ӽO[��g�y����:�?������v^̋9��  u
�O�9\�Yuf76rAC�ڒ,ڇr��G�x�/��-�b���7�~��N�:��⾸����y�|w��}L�����~�4x�slڰ����Uw��o)�%�aa~fn#��D��`�jC��~ͳe��PMЧ���6��h�b�[�
�xA遽T�.���|����[ݳ���j 	%��5c/�3�B�F��h��|���(n�B�'&�)l6�T��)��	�����@�֚$/ه��ms�1�v���K6;���~���X�fy;���$�2�����.�D�\�-�1��6��M�����b�����ͥɯZ�\�8��$;W�s!PƧ&�԰@K�B��V��o-�hs��d�)*��*ږ�B#lL[CW0A��SnA�TIͤB��?�jih����2��2E�ԍ�0��/ޞ{�9�ߎ�D�h0��	���s�М
�j]SvM�z0��b(�/���`A��qNh� T,ED�������sck��2 "�i�ERmeÍ� q�%$���'��T���)���%��@�����V���2�QB�\�׾�UU�.�kX�/c@HRo6������������L�
�H��5��w�t6��ڑ��@���Z�]��m&"�OOMd�7V�n v
�T��1`7sO0��,���j�5:��Ïe�S�2|.�1p���y����j0��Ӌ�nh����2��lH��^��,��}anQ�h�=RQ�E(��$��s HH�D>��p=J+E�� ��}�,�4¥���d'ٌ�m�(0a��sx���{��9=/����ۯ!s4����>�B����vN�~6(3SmAR���F �\��I�
�3ɐ|��Vmdڇ�$f��QӔ�L�x��B�'�8l�g���~�0��H������yܴ6]�O!��w��,ޖN`E-���g�X0��EL���|�d�zE��*	��b 
�8�YЇ]mA���:2���Y��K�[[&���B+ja�s��S�h�3�D�BD��"a�m�!�s3���_��[�cat�!L�|��ݜ_
���VUe��8�;	�ZHJ����k�Y�D��\���<
�/j��Di#��g�u �G�{��i!z1�6lR���̼a�&���h����?���� �9�y�n_Q�@�e1����������|�o�o�:~����*�/=l�!S��]��a��,Q��@��u�k�ؕ��TJ��4Y''${���a�oA% �=�y�'E�oܰ�K�@������� ��I])n�J���σ�YL��U�W��K]�����mF#5h��/{(�T6�_��%����������(��n��|�OQ��|-&LGg) ߋ�^��{�0�I����F����2N<P[^�u�:-^��DOC��SYY���Eܬ �f���vkL3�R�.t�Y�-m>���UϠ$�&5�W�]C��N1���ayƝ͞	P4 ڧe�M!��+����+s���T�B��zXl�BE.��b�u��������y5�n%�ِ�eV֒lU�m���~L�+�YM���Rmũ�6�63)?f�r��chIF�Y��Z�{�e)(]=Q!`ϰ��Q�Gڬ��4{1�[��j{W�z-cë,ԫ�_h�'�>*oj��I0�l��J�'�k�U��Q�,Ь����X?���}%�>�$��"���	�lS�M?���$Yl�h���0+�C����&�k���mʅ(��dm��a&$�#`��0�.���y�}y�o�j�,C�p��Rc2��.��DT���X�@���}��+����J��>����{[��k��t0:'94r�I���5��#U1��Z~i3 �B;��V"������G8�P��`�j��rV��z�%�nI)ʣĴ��6�ߜ�R��ٜ,n�&Yx`�~m��fGaH�B��s�uc�QIL�L7�T��桗�2��G+HW#׊�lz5��D^�/d�?� :W6�>�8Z���rV]��F<o&���K-�\��T�fnk\�8��U�֍-�Mp��&�L�`bi�i�[�F��Zr!]�R������ �P>̰k�N�w�mndl�}��u�5d\	�!��y�`#S�E��&$,y��a*��[�aSTM;�:��tV<0��8�V�H�^ �z�w8񁾝4Z�=oZ&6��Im����n(�O�&*��m�&����͠�Ӝ�$��.���>2S�g]Λ�'�Lx���o�r��!^��~T{��L�6.Q+g�P�L������4�1ɥP���Ɏ����v��3�tdt�|ͫ/���� !
0�h&Th�C�B��9��Ҙ���ۋ�.�
�`�ೀS`�ɴ��D�N�Ѡ N>�L?S�J>o6�ˬ��j>6�o��@�$ ?��T��xs���,�0�dp<���ĭ�XCn����nn��V�}�S��1���F���f_�E9l��Ey��$��N��'v���m�՘��Jt�Ƀ���f	S������D�#��*�ծ�q_)�֙,K-�"
OU���h^k���< ���Z����C=�=.)����Ƚ�Y�iiꂦ
��I�Rh) �j����Px�R�%׵����>��sQ�`6�/��6��	 ���S!ܿ�ۄ�Z�P�a�� O��F?�b�VF��0��[�*����R6*MC�^�Z�K��dqൔ;�P\��DS5��x�BP�l\���2�ɊC��*w���I�Z�7�����_i��ګ.w��YV
n��2�U�(��4��4��. ��aS(ʸ<�8y��ǎz���IHD��p\���uhc��a��o}��ܓO<�:�5�i�A������
cb����c5m�jc(����OC��Pn���a|�S!�0�Ȇj�gPcUmئ\�1������3��*���g�(1%e�����$e	!�a�ϗ�̴�dl"?V٫��lj]@��Z5���zF�TxC�a�oQ�ek
���3`�Kk��~`�KM�����	�m6�e~��4ɀ�5&��s�͑��Z���3���3h-��;,c�E0��)����߄���������\̔0(�Z�*�p�yU#t�1���a���Ǿ�y��v��V����3��/o�g$L�2g�JЁ�!e$�;o�}SV��aj&3������)¤�m���e��f�C��#s~H)7�$�&�T2�b�φ%2�����D��滊�Y;-�U�J���`��.��@��b>z5ޥ��$�8ǋ�w;�\^ ��v_��.7�_zeHT�ȳ9����&�U!<��W8�ݾ}��p�cі@���g�=�1�Zn�_<��L�if�&��
\���`��(����~�񯻷��-�~������Q�ϋ��If���an�yp��w��a"�u;v*� ��h�7�b�By#�ka�<,R����ח(��?�9m��'¢4nA�H6����-�c&��?�;����f�/�YSF��`�.�6�A�s��B	_�i���^��� �JTv��	}������ �DD� /_�䵰�pp�������1��c�4f�w����O��O�����n�޽Y�_�����?�SE�d���(,����4�e�s�Q��Xk���l�N���g���wQ��w�K>wA��>�i�	�
TmJ4�i���L�Q[HO��\P��[��(��_������Oi��Y�F�I:7\��r���h(���X@�I}kk�Y�l��>l�_0��3�d0|&�!""�G�g����h��z��ɧ���?���#���.%�N�YP�l���(#��ѭ�>m��t��t���R���W~X1���<l�M%h_�����O�����"B�#���G����7~��O}�SZ�l�lK�(Pʘfl�\s����o��.�2"�N���ns׌�k��  ��l�P���5�N������krʏ?<��Z/��Үa>"?�{A�?��)t^�\;�`~����p${T�2 B�t���I�6'5�y	�	X�*�Ġ:v0�h�|贳)����j�K��}��E�\���im��@����ϩ$���?�����^(���=�Kiď�@BI�U����}�������Rˤ�+1���ߟ�%i�p�β�w_�rX�~�g�}�C�+�I,"��T0�C=�0��#��?n�{�q�'O�l���a����`�>��Mg��Guuk�4�����q�Y���F!�3�&�����BF����n�;��
�G��13ɰSoٻO��_���H�W}��,�C}��]�aA�z�>�3�U��X���]#*��_��k��)w!�Hv����N]ٿ{��9y(5l,��Tz����>�����~O���ހ<%f���H(��D�o��D�}	�f�h�ae�OQ�!*hB�@�����h;��TefJ`��Ofk�b��9���/%"E�z��H%E�k`\��zp�Z�'����;��~�~��>��GQ˪X O�F���n����# oS*�	�ʪV3��~���vw�VМ�9�jH��两4[�i��7���T�̘T�RLn(dT�cZ>���>rKG����T|�I����>̣v�� mS�n�ڠ ���B<���W[��=�j�ٌ������y�[n����'���/�V������l2|4L���P� ��F��=?y��	˄��LO;F�w�~�p�������PQ(ߺE�%�{�?�v��xf��q��j�C����������}@���[^��w�B��Pt��Z��/����$&���?�l�!	�Ǧ��7��~��o��o�i~�%r�p���|�	ffଦt-g�,w�5�V��8��"�a��
8��Ki
E!�=�D+�n_-d�#��/�<�����o|�7L1H�L��E��Ԇ!�aϝm9��5($R�Sg���q�nc�"����CjA˱��������_u������y���RQ1z�۱}G����_����o��otӸN�/?w��d�J�"I~^bC����Dp��5�Ƣ���w)4�؍ƫ�ηL�G:�K�_,8�V����_����Q�eŹm��)�������G�⑇�^Ԥ��D6�!	�'6�Vmŷ[����	�c��TDA�j��F�����>'&����<��o/#�[&�T�-i�wA
T���ג}Fz�Fg�&���(h+�׹'r�dX�mSju\u��^��#RW�b㢁񽳉5�{���>�o~���2@��4��Q�c�/��u�g�c�����e(����(�F��BM���(�ᙟ����9���r��I66:�>�e�}�)�]��{嵍Imc�zh����wev��B a%����:I��>���&/�.anذ�#?��z���h�>`O9�LiF���&����2&3��Z��:iҬ��	������v�kŠ]���������M�����.�:�����a�qq�"��/jd���R��G(�H͛O�2H.���Rya���	�e�ȼ"�<~nY7"ݴq��ɟ�I�Д�槕����y�G���t���?�a���aXIPԈZ<�<a��ܗ&�D*��O��\��~ӛ�~�(�ζ�3���OPpC���E�U*^8U����a/�zK��W�a�B�����%@�\�H�ZO�DK�0��bJ'#��森�{����D˸�d��n!�dv�&ZE�;���KZ=���u
�oK}T���Ǐ�MM�'�"�"�NBL�t7�5[���r˞\�2���H�I��
�����y��fC����G�RE�Z�oЙs7��A�`f�$�����^��[ϵ��X^��(��{o�q�I�:����=a���p*��N%�s�����R���L�;�y;��a�CG^p��`��>�����s�=�Vc���A�y�ۿ_�W�������'?��HV�Rt/���:�4�is�)L�h3q��c�i�� IL�xo��)Z�R���7�VU�[ĕp�pT&�TI���&}��&c�I��H ��C���|B��n�Q�G=�S|	��MY����(��¼Bӱ��O(�C��}#b�h"̫���f�����Z���"j�.�r�,fqO��������C8�0�@���������� ��0³:S��kQ�D��9u����������~Kg����h�[�/I��˛ױ|m���j VB�˭(W�m��.�6n��sLٗz��^T,e����+a��d}R?s�w��/_-�sN�.�+��]�pη�RWFy�<�[��u��,$�&��4<x��A��^�B걳f��/^������3m���˾W���0\\0g,tK�����=jk/#�dr�"[HU�������������cȗ���}!Ợ���?����wk�y.9����š���b�*��ѣ���'k����?�O*x�%k�m��\i����y�EPX�Ü��`�j&�d��Aq��u���1�������r�0	��G��i-+�q�wƳb��p�SZF Q?��w�}��N��x<�MKڮ<0�~�Pq���Q���i͹h�&�_me-�P��u4�&6�4��춭�j.&k�H��c�;�	�i6>U�u��0&��'������W<�*��3`�a�}S�G��j3���P�R��e� R��3��s���������#�ܧ��3n�5�w2sĽR!��r�bw��O��g&8�@TI���+/[�9�kL2��B٪��g�,�l�y%��`�w�[ǖ/)��POg�_m�/�J��8�����_��_��&�Q�� �0�rփ�?:>2��]�R�}��˦b�A�i�S�����E�N�8!f-�/�2p6D/4':�8;w����%�W~�{ ��a�@�����|��|�L1��e�T=�h]�܃�J�&5��O�܃>��@�˂|�e���.e/�L�hѤK_�-�z�6q.Lp�`�S��� ��Y����s#@���ݏYs�f�Vc��1|�)�H�qY���%1�|�i�J7ݴG;"�!;�� S�/�>��>�����X0��R�/4S��f�������J(� (��9pa�ة26�L��'~��f�O|�:��ˮ�n�Ce��l��5S�D��&���95���?����{��r_��ܺu�]9.��o��4���֨�ڨ?�^j�f,�`���)�Km�1���UEF��}��a�XC��[QG|��H��o�׵Bxn^�4�0�N�9�L�(��l��O�i�8�/���Y�S�)�k�<�{�����]w�y�v3jNɑ�54�7
�5%�O1�!0�0=ݺ`/{��?D�KC��X-�7P��w����g?����ж�H_��f~ɾ����ǭu10v*(��
�i��kk�Z������>�:�k��z`���կ���dq���1�����F|���1="W��-���u���̹#�_��1��Ѩf���u�y���em������ul�$���w��׉v��/|����7����i�>�}В����~�i?�a�b���t��+�Gm_��>tD�# ���[͖��됿�c#nJ3�s>YV��Px���������C��w���#��5������5�0a^<rL�fvf^�ueM�#l��##c�����������r4!�Ry���J��L����A��f�ss�R�;�d׻C��}��O���z��O}�����0���2v��pD�7�١k�5?�YϯtD�Uj���:ld�hpp���5.�׳�9��J��%?3�H���u៕�D�G��(����^�Sk�tJ����B�+h�Ŗ�=���^_W'��^S���g�9��۷7"$�Z��֭��'�p�YG�k��R?��B�7����o�ڃ$������c�1�3���egWXtD`�$A��eI�R��R�R����OB�l�!���`�
UhH��-1�R
`@�ed�c�g��g�qO��;�����3�=���3�V��Lw߾������xM�?VYq���a'�0'to���	&�aD�Ji�!5�fB��"�) T.C%s�]��F���0�i�m��S��cS���{*r�)&U~�2q]�uiPh�4��9btOHO`B�!*!���=~,�y��;Vm(�n�W�n�$9|����>J�zXؘ�{��=.���o�:@� ��F���]k��'���y�N���	�I�}��%Ԣ�g�",�V}�0&	`;)<��@�&�����!t:s�ϊC�������	�0b�d/�rH���P:���6�A;p�/F�����4��y�D����������&㡡k�Z-�KS���:>|P�{�����r�b������x����@�a���yf�fѰN�ҽ&��"�n�d���_�mz���D�x�9w*�G�,�Eq]
Q���I�O �*�*��+5�㡆/��-�����#i ���(�<��T�?ݸ�G�}�J~\�YtL�����n=��C�+�o�0�Z2}�b�1�������m�z�Bc�4[����G��I�H��<PT�����p�6n������R�MC��A԰�!�i�<��in	O$��¡����co�x�!���E�6!���?��ω���'�[�8��� e�q�`E@��8y�-�o�-���z�V��X=����D)�R���\�����|>̒aNvd!8��{��R��}��/2��j��}�=~�,�ӓ��[TLH�a�#�g$l\d�ӎ����nC�C^r�%����wR�|#3���/���I�W��b����`��u�q�K��Y.�C2�'S�L��0@|<�K�{�;�/,�(��K�ju��_�i�!�5g�);n�X����(��I�8ݚ4�]����Dܺg��ԧ>E}H�q,A�n�` ������m��&�z�)�m���G��d<��K�[1L+󉚾-~�K	q��*�@���\MAlj{��If^7�����Mg0�CZ-�<�a�~�yc��`�H���r�-�����;�y�É�v����g&'��o~�AK�O�Gi8���`�+ƻ_����@ Z$r�f� U0mo@� 7!���?�"B6]w ���q8�V  ���I@1����&�l�0��H~�^���CݫtB� �Ѹ���mr׮]��ũj� 6�O<%����}/�O��)r�e��aꠤ��G(Og��4#�Q��F�z�(kdƣ���V�=�:�!����bj���	7K6�����mZ~N�<����?�1���e��K/u�uFA4Еz�o��B��|	��� �T\�^W&�ɇ���c��,��:���Ѵ4�?@&��7�Exɠ��)�s�C�h/l����F�����繨��yn�4H�2E?�я�}/�	�s����Z�A�J���B}Mh�W��k]�Y�����[	'M@�0��A��Ќ3��I�����q�$�Z��N˺w�`Ox�h[$�/��S6=:+����,��ؾ$7ŕ��܋�k֒zB@�^��	���}������D��5�\#?������Z#�=���a�:�����[~厯��w��a�1��#�5�>Рr����{$�{��>~�ؾ�"���ļ����<a	=�2�#\��M�+)[�M��K/�\�~���:�C�r뮽^T�b`�pM����V6�)�;``�l�:�Lߌ��zA��7��T頾���Qq�w�q�F�Q���-�i���059<��L%l6Yt�����nr,��tM��ICy,����|���A`.H$���g̓�7��g�Y#N����*����7M)9��$O�mwm8���YR2����.�LuϿ�#���oɏ��Ǩ�x����2o
js���G���GݍbQ0O�E��ݙ6�1q�)W��<�x����
e2��(�bA�� a!w�R��w��x�'�ʜ��Ӡ�҆�2�mUOC�kߤ-��i���G)�Y������}Z/h$|Q�H���41	:�;��p��!��\ޫ�$3U9��2l��j�3�'��uƒ��-������M��g�kh� �����u��a�
;n����j��3��晧���hl�Q%�!Y�������\�j� U���sӍiuq��z�6$��~�[��ƃ��Y+�ҖZe��F�ϳ�=K�C?��ư��*I0���i�9��������??����s6��6��y�z=�rIO� �	�S�|*m4�N�Vo��)m��b�~����x͡�S���ZA�pg��j�]��wh6�9���lj5���0�6����6õ����N�Q5(/@f����>4�d)L�2&6t\?�y�p9N�ﵙ����fhkf;�7���{фA�N:�hG�9��s�#���Wdq[�R!1QX���_�������}b玝�
�`zz*�90&lx`h����[�t.uxhƠʷ"lB�CX_��kn������Jim�ҥl6�y
���?�Kd�y����?F�I� |`�2�7g�>�n��Qf�f�)�`*��0��x\#O�w��k|0D����v�7Ȧvl,#���d:%�b��u����;��s�~�L�ŀU�̠6,���&�.M������J&�4��x8.�k��p(��Y,ZH�$��!�����s���L?g��2{�� �	�����_�׏D�ۨf>[i7��~�i
R@��]��Dm4��9�L{z 9�2tV�rs��ъA��l�j�DscOE��@,"Nvș�-���-;�,L���טh�l�����4�<�%�چ����v�u�˟s����5aF�����b3cR ��fd��[�̖�?�� ��n�����{�F[3 �i6O1k���b�z���%7(˯���c�o�x=D���*U�O���L*#~�z\~��g�yZ�V�;�X|h1�)i�7;�PF3p,�����4������I���-�#qq1b�am�V�EEX3���ٚZ�a��W�w�$R#?bB��)��y�3IR3!-H$�5��T"��K����+=�X������(��`(gc�E�w�q�bH���c��EW��h�2�ڷz�å�;��9��}-�h��ܬ��u-��z��}Ɣ��p?��k��Z�6�C����k��5��PXw�-E�@m��귉�X�Ȇ��N�ߖ"9���N�Jk`D8�.��q�͜˚�c�MP�`LP��e����V���_1���%�Ѽ�~�q�c&�`�c�Y��ơ{�뷺�Ř(~��k�^ "�0��5Hwښ/��m2��F�©��C�t�� '�4�gAr�������* Z- I"ሠ=NfR��&˭d`���64��E?��u#(�f�j�D�5"������@�T;��Ů��%&�ri�=0�s1�)�<}���P<j����w�#?<'{ ߚ�F�nDE��b�oZ��T�ޫ�����1%0�d�9C2�r*����[���Ry���7�0K�ڄV7]��'h�__�n�D�o���^�m9��c$�����y���(s�`<k4�	rN��W{��fU\Sb�J\F%l�C�*y���^�Oe>F 0�����\��kF�^��9�������a<z)�M�(�q	��{6�Ʊ���x�m�7���S�\����G�i\���b���3ωI�,�`�ɉ9<uet�E4�I�^�vl寰�Lm�xݑ�,��M��V�
�����	��di,D��v���T�0L4�Y8L�w69Xq�0�U#<W�Bq���C'��)D|':�5�m� 
�J���P�?_,'*aC�3�����&>.#����%�v�W�E����� 3ڢ]"�U��El�1|=��w{<�$�%� @��=!$����W��=�q�i���o\�Om�(��rh��L���.�ɠ�e���(�a��_��ƿ�x_���H&�'L%&��K��d� W(\�%�]�P��-G�%*��/Ď��uS�O"h�q����p�04ք�48W���a��r	���D��lihԛ� �̿��pp<��M��K��$��������sZ�<�m�ɔ�h�LH[d�!L9��I^Zk�oZ�Yӥ^<��m�p�����/�t�$?�ghr�I`#��}4-��?o�����r�D�8��ؤ(Δ��0�!fG��	y$N����tV\��Tű}�vƔ�2�	(��D$?�+��K�J��K��n>Z�4�\P���������sjj:��A������n'H��'���Ͳil5&&��M�ךَ2�[�Aش�$�]������LV'�0m�`T�b�-�����;�E.��S\����?Q ����~��x����3�!�L�e˖����I��q������矧�׽�:�7occ��C�E��#�<Bh������ë/���(�Mf�^v����7n"����d:CI^ɉ`����Zu�#j��LJ�z^��E`��"l5,~A�Pӌ���o��ؿQ�\OĿ����ew:�(�7
3��A��D"+�up���I�o�0�T�'�gB�(�9�5��j?Cg�m ۄbaNZj)�
z|��l����R��#�tljlt���P�����$i��PCk���Z� (�4WA�ࡾ㋯���n ���s��㚹��}��c���(�K�p�Q�k�.�B(����:�E34�D8�Ye�����%���^3��z�8���:Z�$D���賵�5z���}L���\ f�\y�◿|"��M@c�L���� F�>J0�79��f���g��qy��nB�/�V�M��QZ��b��I�焷��I]������u�H�`M������ABp�ؐ��v�hæ1Ҟ�_<�?0QR�]1���7�A�L���ؽ{�����||���gz?�`#���Z4h}����f��&LW����_p�#��z+��`���EG)��Oa�a�r�-��@7��P&�@6b��u��D	,��h�d�T��F�O&��x�<[X��W��{''��P��)k&<-E�����8�V�s�F������rn��v��O��P����t0�HV�n'�`O�{�{ ��y�h�i��1&[��	A���d����e�@�֫���U�=����gxN��T��	fX����#�M�n�Z�g�gi����/t���/GGG����E{l{��8dN9��fK$�S�[�$(���GG���Ãz�-�\��ɩ�/��B*
�$A]z�\��s=�@�㮝�N'���ڂ2�֍~��]�袋��4��Ø
��8��dmNN��V�^�	�43�l3�0$�Q���܊Y���m5Z��i~K�d�{ОJ�*����#�|��a�o,�JM��{��CC�;��I=KƵ �D��C@�jH�&�K��)�z�W+��*y���
K���&\�iJ����+.O��`2` қ߼=xo�ap\Hp�͘��?ycA2�{q®c�oV�A65��P��
�{���g�[rr�r웯6O�>���r}�u׶�y,R�#���z`�<�LHҡ�A
eCs�p��~ ��Q�Uox���UW]�(F}�h��yB�C��'��Vh.����&�g߇�F��>F�eb��[io}��Ӈ��S��ЈA�裉 y_��5\*�I�X�$��:x!L1k/�����T�*4G������Ż�z7��)ðd����<e;�߼�8x�e��ӄ�$����m����:�@0����p�O(u�cQݻT"�Y(���#]�`Z��#��ۿ,>��^ n,�	��������&Y��;?�Pz��\ij����>(���U��c*�k��M�E:N`e�MݘDo<n4y�/1Oߧ1<�/}�K#M�aafs7#3��0lr*����N�0wڿ�c���<}L��uF��̢�Ѣ�<^�>jk B:���gQ�T���Z��K���Ɲ�2a�C���d(l^m�b�nq|h�0�s)�4�6���o;O��&6���s��TB�f�6e`c�}��B=$$<L<{���M��7ǌ�Y�&��5��_��x�;��@�q4fw\��f�M�q�}���%�Dm��1ej<������PVd��:��3D�se��20���J�M�88���u@O�k|�<��m&����9(�������}0m��,/���;gC,�<OXpx���R�cK�6�9Ue�$�#%�s}GD*3*Eo�����M�t�#u$�4?�,�\e���f��K.�H�>j�����7C�6����0ܙ�E��XD�i�����^<��)^�wBz�)��&.��(�R�u>?�B�o��`���g�~o���P�U��D�ׯW� ӘWL���rc�{�]P���L��>�*�`;��%���o�ؓ�L`��y�$t���v5OB��ֺ�P۲e�#�Dm��iثb�L�O�1���)���)Z	��8~��Ț��
ʬ-��z���|�zڳ�"����$:"I-�9�P��l� �8��x6�u��m��ƂB���]�r�����mO4�6��M�+!DD��C�!M��yhUy��21r	��Ix>
*/vY>S���4�߭i����!,%dU�L��KhļҚ!�8�`J!�2Nec���{u���Poh����0��_��R�w�Q8,' n@쪹�3������ϱ���:�ǥ���������q�.%��`����Dɥ�.`��o����mb��>̩YPٔ�>g��������:V�Rͷ����^	G,��{0����V�ϓ��Q`h�8��l�k�t�#��#�� yoQm�T��  ��o��g&nU=刪�r�H@��#�����F<�,��T��H@��c�)9W	��lWr9��0�.SK�i]��X?C-c;�T!�lµCkı#�)s�j�X�cǎχpg�f��NW(g�י�)goG"/f��y7x�цT'���Q$J����!!'��+dc$w�wLaa�����\��J�Q$0�"��kb"uχ���@Q�9,���`�4�#;v=��a�y��Pi���!�	�����A��{q�R��N!��¹���yju<����Ԉg
a-��AR-20Y�5�z6�w��@��O*�cnVO�C��p�=���3í^_��;�6�	��I��Èȓ=3.�r(�>��y��R�{�0�Zu<�p&`OC�HQ��ȸ�[#VUK��� Y�_��.�-kUJ��l��6�er�,q諺RG�Q<�I�G��5|��ٙ=c��dj��]�?R[�טTssd��4�u�R�.��{�����юO�	��K�t|���[_~/�s��"�5}.b�*��9�(�X�;�A�_�~.XE�Z峸F�L�$
Lu��"�e���N���A��1}�b�!BFP?��^O�fES(f�5a��@Z�@��QP��U��ϻ�����G`���[Z�>L+
��=�Y��&IIrd3�c��
"�IR_R��Vb��@q��0>����C�$�䙽�O$�!8�T8�{pŬ���1���f1�D����a�q�,&�u�H=dp��
���2�]3SeQ�T	/��T�]e�%ɔ��Y/����'N�X��k.�Z@� �h��Yu�4^��s�i���(r���_3\����$��\oFK?�n���t�4��6�
M$�B9[�f��(���ޛ��#�D�F�,Rz�\.QY2��
5��.�ih��x�~P�����[�p��%��F1Ԗ���Ng	x�A���9rru�q]��c%.��g0!}�6xtHf2)���ݙ��I������t�Zm\x�D�f�M=u�aK�)�eeQ��ăf$0�:��t��o��sZø
�e�N�a&�@#7:A�|�BH����)��`ʳ��5�ݞ��c�������k{�0>!���х�(D�؉ �F'&�І�ieh��o�PE:�W֗#:"ʥ���\��:.1��N- �2ו?�G��N���R��>��&��>����^7j�r� @�#�9�$M����
��;]�2LV�Ә�^%P���D����E�_�Gt�;#��3���(P�<`)2�� x.֢G�i��ƭ��
�q�����Q:����d�P?�
(_!�&ݢ6W��V��D� _���k��>5}�I�Q|f��d#V3�l���Kб��?��j����W�Z��t��L������zѣJ�ʏ����7��ap�Pz�4u���"�J��`:!�-��)&!�I!t���<��/�R�ާ=)!\^��Y_��**s̥�1��Vj�S|]�O�c�y����P�ԃ`T����������d���B�v&h��M»W�(µ�R�!�fD��>�#/�	m瞫�Px&�/üy��3����C�̸D�%"��@�R��U�V�|�L\ǌA�^$�{�
����NgD>ׯܷ��x�u��P?0�M	� /�]���]?L�n�8��.=][&bP�PA�m�3������q�S��.�'g0�N��|Rư�W|�)k�# @<�D�J��m��0��jPr��O�J�}��x��!��~dm4���N�2�b���P-O���:4/1�=��\6��O����'���-c�ءWE6?�&!f�N�ɩ�J�Y)=�$2N $�?�CcE`��<x
�"���/C^+�b�zG�+=#��|���_�� ��q�����QqbrRd�fb�$��ŽJ����ߦ�ܜ�SR��L8��+쮞$r�����d��M��c�mo�.�ʂ��|M���A<�,���b��ukx֨�l����ex6�]���˫���|���1V�@�ض��,~��_�C���ѵC��?p��Hx9177�I���PA���,�Y�I�fg�;���~3,�Q677��3�#�\�v��qm�F< ����<F≯0@~+��A�~�Y�?�ay�׾,^:0+��;�,�qَ?LM���� H�b�Í�pbw9��&�&��y����o��k2x�*-�0��8;KC�`�"�y4�qL-�
b`�%�liZl��B�/��+����Wk�������i����_�췼6�1o��ab��;�,+S�&���UߥS2���)�~�84����e3���${!�\�Au6a,�3�����}vb��r�S�.�G�)͹9r�bP�.�_*2������n�:���g>��Ʉk"5�8>yB�f��_&�Y�.Ȳ�+*�9ED~F�����f�Ί�a0���'Perَ�_ܶm��_>�(��ǌ�?��j*T�jo:I�Ӳ���a+�K`�33;/���\ALK�^�~�i�G�L�&L�53L��a>�'��z����F���Q����B�Q����<�I��� �o'��O���t&S:��隿���*�Jf����$6Y��ץ��3�O��p���'K�e_g��<B�X:6�h�ڥ�i��PݭM����w�]��?�Ƕ(�w�2ɲE���ݕ�mN�Z�g|�1��M[��n�G�aq1f���:-�ﰘ���L��2�R'��?M.��b��DJl9o��&j�-�/�׏��G��H��i�f��s�i�6�I�0�Nl�Q��=�� 9f�pb�������4��k�h��*uJ�:�Q�T��eՍΊ͛/�/����_���	�O_�f�g65�f�Mk���4N���p�_���s%��z$�ύ3E�c�V��|D.Y�XKhpI�)�3�7�J�=x5���G�egqy?Ȋ���B��&��cg����s�hdig    IEND�B`�PK   sRWZ`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   sRWZ� `�5&  0&  /   images/e181a1ff-876a-43d9-9539-3671c727f4f4.png0&�ىPNG

   IHDR   d   '   vLz�   	pHYs       O%��  %�IDATx�ezp]�y�9��w_� QH�{�XDR,�%�*�R9�S��{3���d��ڙ��Ėl��Ҥ$ZES�H��� QI���������I��˙G����s���_9�mۨta��b�ڛ<2V44f�����XH��$�pѰ�kc��/Cj��8,&d��8�**�I���my(�p���$� aG�3�h�����m�B�NVul��C���B��ӦAb�B$�4/C�U��(lh^ʡH*�Z��C�z˨��C� ��^��HU-��1!+�i�Fb��pPF�{,��l	��fIw�O�9�c�B�dM�;�C$�Y�j�<m����w�E
���e�Z��X��SO�{?;�q�d�@������}��3g�'06]��O�T�^��L^�0�+�w<�кS7�q����E�7_����{��]CQ��7���o�h,��['�\&�o=��uiÑ3�\�� mCC�Ϟ� �<~/^����}�߾�Z�п�������?S
�q��	�A�x`�_=��L"��wN��?���-{Z}�FϛWT�Z[�}�'<4�G/]��H�����o[�����'E5ę�y�5��G.^;|�Ǳ�-M����~���Х�I��5u?����53��w�����B�0��f�:���h}[��G6�n��ȃ,��9={cX��'�oܼi�eY8?�[�\{`���E�M>v�,�w�X��#	����		��{vnٴr��t���������Gl�=w�OӔG7l}b�V�����GN�����}h劶ŵ�]���ٴ��'w��ӊ��}v���L��k��3�j���<���������F�h�صa���e�E�+�0$���5;��]�/^��}�stɲ����	��؛�}��޲���;]��._TW_Sk9V}8��ڕT,�Y���Y���FN��$��bScq>�\��-��������Ʀ��H<C �LfG�^_�V�pZ�XK���RYQ1���C�� :Y0��⍎���abݢ�c�
�:��5]VL&eK�c�TW�ka�`���uu��ۻc�4���ᙞ��5U�n�:&	r`6�#���L��q3���wG�~��힜�<$}�J��[�F"Ꭱ!Y���^�nY^?>�J�HOM�]�վu���C���	Ӻ����S��'LluO�E_�g�z�����ĭyt�w2;�?��{�o�G��������(���������A��O����cՑ�i�66N����������<&9�a:��t��2iY'h�w��?�ћ����H�k"g2�~�c�hlf&A"֤��S�nvD�y�h�6����εOE�C��W���'������t�>��]ꝼ~�g��-��:�:e#B���a�?���/��	�ri3��ʪ����?}Ya���(&h��M#��Λ���-Y��of�kx��r �1Rr��7��T����*occ��c���8C�x�l��u]�ַ�ۅ��+�\����sɦ���h<�m+ey��A"3�5�.�]S1���fB��*�l��M묥�6V�{��;�~���?���\���D�R��[�1b�?���r୓7)ª
�8�//��L��p"�y�>!��'�]�VԴpmu�iX�|qq]dIu�i���f�\dz6�ʋ�wu��VUI�|M��w�3UuU�xv��5+����U+�-tg(v�ohM�?�^I�yxu�2a"%Ӣvwj��qMuu�B�e�B���i���h:'O�ss�����+��niYE�lt��o(��+���Ics�`��|<�a$g�����L|4��DK�rS9�W��Ŕb�>�e�9I���)�c,�3�s3��{�/Z��Ide�d�f�l'�d؄d�$�����F�&x���� ��Pp>��>��\}�?K��B^A�g�᱉���)��`�)/Gg��՜e�;1Sعqɼ��Ԇ�%�ض�e�6I8��3��$I9��h�"٨-���l`��Gn��z��|ms�����b(�@�U����E�\U.�����ɬ2t��ȧݶzx�80=힗�12U]o�� �����1�!�hi�;��񕎄�id6I��3�#&�!�$���|A�R�m����O�I8v����`�Oc�"	�!(��������YΪ���KQ��_zqWT�������6���`τJ�I폊E8��:��7h*T�0~{�� ���0�ʁZ�p+��m�4��!Y�ab����e8�>�q�O�$�n��z2�l[^��v�L���=54�1���-��J����Ȥ�>k]�2-{ix��,K�0a�*�39�� R�<�$#�w(�a��Ќc���poL�e�%r[F2M�!-�2�(�\���^��r(�Y�~�+�y��]����D�T-Ͽ��ZY�hN�޺3G��(vWȲ��U�V���y���&g,�6,� l�"-�^�%��Mf�_"�9�h��J((�O�>"����Є�W�\��"�ʖ��:7?��ݛWׯ[���p���'���7>�5�Q��-�FXt�Ca�v����@�ؽ����"��&E�m= �5՞r���Hr<g��a9�� �t��Ŗ;�i)i��xi��yp���n������遮A���%فѹ�����	M��;ɬ�zU�7I��i���bQi����O&��|6��{�2�8l��xJ�m E؆�uv��]�c����4 �\�EB�$߳�nO��'������o��z���8t���%Kll;t�^���1�hY	,�"���j����b^5a��ML�]d���_"	�����%$T� �BQ$��C͡P #��}��/p���B	�5��ѬėGX���stV%�((�iF���i��p���e�E���l>�gY^������Qk��}�Ժ�  y����m���S��B���#l��r��@.��,v?���J��l����#;�_��g���W��N����4A ����8�L6S�z�O�?t�{� g$"�\�r�d����y`H�!,D�yY�>�c2)	�n�:�h�� �b9��6d�A���@	���2!b e����?@s�T��p��h�H�-���b�D*oa��tM�
�$�@�A��,o+-z�mp3rR��tg�G�`8�/؄�b�J��ܮ2 8G"��KFg�mXr�����r�F2��U��(���q˔$�����C&�s��#�k����$���0��� 9:bx��5)��uQ�1Ǻ�F����ʖ47rFjIY��c�D�hjm��MGh�"���0U�o�2���lBٴ��1��
��-A�B8���K�7����R�����;7o��N�۝�T�P1����X� NrddxŊ��ڠ` Up� !c�ӎ�cƂ{�4�a�[%�s�^�i<�KR��͹�Sݵa����\�6Ґ}��ӊ�0@��i�������m��<Ǘ�C���ƺ�۳29D`0���t�!ؓa�#ޝ-���&A�!� ���R��7�ޚ��'v�[d8��JkV?���}e��K�6�Z�L�z��������<��N��(���q���~6�@����G>����V��'.���/��Ҳ��!�9��m��&�������ݻ�jk�\��2/\���'=��U�k99�!-ҡ(�e]��v�3 pͱ�l<YV�К��6,i���xx냇~�I�p/��`d�$���b���nܼ��ڲs�#��|�侽�Sq)��E�"(�eM|(=���dR�����f'l�L�b0��p8кb	�5����gg�!x�R����?>�^Y��٩�8 ������ �P2S���"A���;���ݤHb"/B��rҽ��Ɔ�DN�U�Z�BXƪիuMmjjz��'�[��]\!Ĳl(��sVNA&�4*��K��q�]?KP���<B nRL�x|�@oCS+ږ���A��@ ���_������s3�3�}�ȷ���w�_T[u`���DgB�(�������v��]��U-*���ۆ
s�r���s�'$ǉ �wNs�Ώ�]��aٱ�b���7o�����5���\�$߿v?Y�����2�7���|���ᑬ4��)�$jP/�r�]�sXl�iZk׮iY֦�q057#�eI���Z�"�������a&�؋��'v-��ɩGw�y�}br��=P)(:��R�P�����Da�S��W_?p�qQ��\8���w��HA��L�ϰ��F�B�0$����
?�V�U'h0�A��]Jeb��+�j�g��c�_�P�$1��v&]��޻uC���c�����$v@M0�d���y@���+Wx���_�`= 5t���r\�kX��J�L��^�O��%X"Oy��w��.���ms���ɦ:�rnx��՛�TRU5�t��`S��&�kF�4�-�Ka0���[��ȶ;{G��'T䡙Ɔ�T.���/ h���~I�vҒB0L�W�ꪒޠ�J;��=t�6O����[/6��,H�}���GU��M��tMw�xJ��Ke�� ��iM!}aԅp}Y�|Qʀ�Z�J� �5Qxh������ꪉ��D�eXb*��pEЁ���B��J�#�#�S����+�`��*�%������h��� ��"�`�����׬����#�/�~����]�	R�%EVU�=���h҅ |��f�������ޟO!��^��eʿ<~+��J�ә�A�z��l��8ў��u�`��R��U����g�R��~r��}qq���ܽ}�����?�1�&��n�R՜ҵЉ�6�!�	?���Jz�)P�M������zy`YD@�Ţ�cL�w⣳R)7@b`�t�c% �4	�r��&xA��qgOOΓF�-����(�0S[a�G��k�U���r��\i��3<�d�_!���4���9Ӟ�#�"1�paCs������	����X7���e�e�(�~Y�ف.�t[k� x7,_�PQN���:���J�=/�$i�e����4m�dЂ(����0���&���gΜ9) ��@�����d�/x.���EUQ4 1`��Ȼ��jX��Wwe�V��Y�@d���0��z�4`��܉��s�Qxd����9
+K[�]�;����ɕM�P�|!o<v���7��VW���l��T����NvB@x�j��j���{yAQ�cW�wK������4�* ޞ���@�^��,<� �����	Y:�P�I4M ����i�(i#D��镲�ڪlCij^�������,d:������@r&�X,�E�
bC3w�ڥ��G������nǆ��si��X@�qM0v�LP7�.`Y6l6�X�ú����6ז�M%	d�[�ܲ��G2��(����w^�۱f�dN��@ۺEݟ��
+�~#N��_|x�S�2Dq�H�v�'� |冀��@7(�5(����/�� � *
��Y�ʄ��fT�,��������ήS�
����l	�ЃC�DM{ ������9��7�[s�FG�j���-F ����V/��M��?�+
fhh���!�0��%�14��#�预a�=EĪ�3�ˏy���5���ݕtc�:��u@�	ӆIj`A,	��G`钉�fJ*�p�� ]�J�n��h��4��7���㉱"��P��ځ4,���s�Ļs��2�Ggo?���۷�ʫ�4���ۣ.#�b�v���G�ů�(��!�����w��]��ռ���s
��Ki�C�T���V@.��3�0EQf8H���a��O(ڴʠ�Y�L��B�J���Z�ё�/)�vδ��y�lUWM���Vx�۶E���:f$zy���n�q\Z�O�LPT�1:6��r,678pY[�޽{i�wa,�ن�S|U ��riQ"Y�D�w�O�z����P�=~�c��&V�u�������_��t6�
�D��
A�7a%��T�T|�+���w|h���|����TKE�P4���t3)*�����d:�+�h�X%,���"�j��~xiy,�U����N\�'Գ��>���q&��l��u��.�i$5e,����M��Ƕ��gw#SO�_��y��v������Ʈ��Rr������)��ݴ�����@�`1�֬jk^���Iu� :1/�=�@FI �PS(�	 �D��`4���~d��+8p�ʵx<�Y h`�b����cǶ���c�Ox�����Ld,�fL�_&!>#SVx���i�@&):����d�Oضm3��Wo��Q��d��C:�2�)�V4]�	V5��j'��鬜Ȁ�s�jmn��@�ؖ�X�"�:O覩ɢMNڒ��$竫��\����|�`Xd8����~Q#	
��D�Y���|b8�+�$��H�-萦K�(�Z���Z�h��5I��i�?��3XS�����:�&(���5}��=9I�m_�n���:�Ʌ<B.�B4�����=�1mC�qk2��z�He&�m��{cj�����
qy>������3�b!~w��Q]E�y�Y���]�za֖�8�/�27q�|�l� X=�?�h!Q����5�Td�X���|��o�����L�^��I� ��$ȇ���q�C��Sq� �+v���%pݖe�$�u��GH��Eʇc���������-�{{�����$��q0�d�R��;֬�|�+T�:�7��LyyH�u�``��
��4,E�%� ʏ���|��U��5Nf��w�}��0{����`��dٱIW�=:kSX���L	&t�v��8�?�3K�3^h��A��5kXde�U�(�P8RU]�I�n?�a%�E��`�?�s/�B������q�c��x6��{f�p���x�Mך�t�L�db��IQ���|����]=u��˖6~������ ���~vdj�������~y�c6R��)om�����cs�,A����D�詬�J����Y,�*��pV��ɜ| �g�$0��	U����, ֡x������qa�`w�Y�.���G^�Ұgcm*!�-�?v��%�R_�\�1��9�}Fd�y�Ȃl!qêU{7��MߛJ�$�,��RZG����J�Π1n��,����37[�����n^��w������"_鹃��n��5��~��'��p1��U��e�]�V�Xz2۴|#��}p���u-�2��-�׼z�bQ!:ǳco��01��I���#��C�&%O��]@z�=n0�aQ
GA��>G�����'�N�|���vL��f�����!M���c7H!n�!Q�gf�^�;6>+x<�(�PN3ܝ#!����e���v9�����R�4G{n��u���_�z�NI�y����w��������#E�4��Օ́h��A�Sie
���xT%��������K��y�e`C��9�rg�E���#�����,�NV�3�:����L����ղ\�LV�cJ'�`����َ���5A��&�ߏ�`PpU�IN�
�D�%���ij����^�Q�g(��E��t������s$iy=4���ۺʐF_�����#�����)��8���l����̍9]���j����yo~Z��Y���?�̎O̝����B� y3SP�����UU�HK�y)	���8>#��\Ѵ�����eao���fZI4ֆ�/�R	��8��L׆ByF���$�JUU��hsY�b�����̼��Ն	��Y����>]��c "�!p�rh�!�WU����-])踻?�n�zMѳ��|�mQH`A�|_,*9YO���ğ}��Dz>����1',k�ػ�gx�s$^ �6������!�0�D�E�!�_>��s�Z���|1�L���/
>2���w�f���|nn~<W��>u�qs[���Y���k���~��M#��Ïܫ�/�Z
�&�"��Ե���Z[
m��|\E����6W/�Rtq"-]�پ~E�%k+˓9��7�ں�K��fj��n�W�d̈́Ч�+�HC�%ݡ5� j8��BeX�6�tkv|z>�(�juu�i����"s,�����sw|�!���	��鄤��mkb:���9.��/8w���H@�^-��4�|�ؙ�ڊ��� �9�5�ܹW�'������pĻ�?�*��
�ffA��O�ͷ�VLO��W?���^�F��d�ȋGO\im��������[����G��󅴁��U�t�W��"0���ڙ�X>�	S˫6��; �[��%UUB��14��1K����u�����3�o�n){rˊ��c�FȾs�{��M�cx�V��qV6Wl\�n**�w��9 ��[W575�N�jԼhp��M+'���+=A��٨���}`�"ݐ��?�e�_�5X(ʑP��c7�l�dS����u��η[��ljjr��}�%����f�E5�ٺv�"Y�����Tnۚ%�7;�q4�H]c�j[kʑa�K�c����6mZ�����"�sɉ��[VJ�v��=����7^صeE[����;��b9� �ZڳdYcU���g�|��������b}}��5���3��<�g�_���<���ߜ��ɿ���� ����ϣ���-���/<��@���Û@�_{���=���w/ԕy��?���n�\�����s������<�
���~�"���WV�5�$5Q���]�;5��/>��p+ZZ_�᯲��7�{��_z�4Dy�k5������%M�M�~��_�7nϚ}�k�jB���{�#���[״�b�_~s�N��M?��K>�oɢ�W~���W�]�'�>�l|���ǟX��m�ACw�Vލe�O���q*?2AR �@��!����$QtP���`/m��łk�0���2��-Ҫm�˒���ˉ�fA<��dA�d���E�&Ez(�*S��@��d`_��DbEK�"��-E�ϒEC4� hIV�2I24�A��90�����B;O�%�/Oed��8�P�r��!�A2,J���%MW
Q�Q�]Ua�h ���O��g>�Y`�1����S�֩�5���bX�������UK��ߛH��ߩ��PX���~������K������|�;������*�>�=�3�_���KYj����uC����kk�yw<&)�=v{��?����[��#-���蟘����&ـ�=��ޛ�Ԕ��ӟ3(�o\�I�fZV�v��~a\������m����E����^ �=q�W�p�C��w�;�f����|���=3���7/���}_aX��}�=2��[�ٞ	�����I���U���Fg�M��a�Cd�	��=Z�rCh���,2��FSw�]	�{v���wF@Y��C���꽗�i�bx���N�D�&(�f��d�2_������t(�}6{~�
A� '�H>|�� ���7�hV���0����Y���!��>E
^��=�[�]��@�M9$�ߘ�ݜ����'�q �8��F��c�!��_�e�{��$�RAYD�������4g"g�h���%�#|�)�d��N��#��eC��j��$.d�    IEND�B`�PK   sRWZ�E����  :�  /   images/e85fedc0-029f-4b1e-9a1b-73b665cc1a4b.png4�P���q�S4H�P�@qB	-

����.�^\ŵ����-�A����6�����ͽ�<��lN�SR�H�K����B +�A���`!GB\I�`II%YII{G�o֦((�q>q"2���b?9	]Y7bsZ�%���Ԫr_rԱ>uf�J�ol�6Q�>h��k�쯱�*�ùT6��@���ӣ�ͣ�k6���7�Q�.��@[x��5r��=�F�:5W^��S""�cc�ǥ�WL�X�B{,�X�3� Ǥ��R��&�{���p�j�9t����l�*sd�4��`G�O"��-PaI�D�ĳv�P��/�:0���@��7�3�$�d@�$�E�X��:�*�_���7�-e�J�LP]X�m�n���X>�vcL^k��R�r���Yx�Lդ��䉗����g6�c��[{���"k��a��\�1�jh+�i�]��<U;s��c�*���a��e�����W�3�|Q�����E���e�������	�38�2�N((\���P���\�'��e��@n��q+w�)*g)-gI;S[gIGS#gӯn��e�4)QPPd?H��/�m�-c�sa�z��t븎��y3���:<$]���ڭ�ne1��ǿ�����|-}��$N`�W/O��-�BmTj`q�_��vY����3"y�����Ʋ��H1�O�i*���cB�WO�YN��������c��P�E,9��8���C=l���?G":U�[m�*�;��:ƒ	����5+K���^c�o���=�^b�ceg��7���T$$뀛&�)�`��A f>�U�oՃFaL��A�p��{X^�+�˘��w\��'�g�)�ޚ�P>�Ӗ���蝤�d�����4
�)�e��n*���O�8�^�wJ*_������"�'���=���!sH����u>�g|	rj���4��3̤�'zfb��)�IX̟���&JZ�����<|~����c c!����!c/'aλ-�����)M�N��HR���y=�"@�h�dD4"�ɯ?�Fg�z$� �l������y/z���D�j�*P@�ϯh�<�#5ى=_����D����dA�����)'%CF��{�w�Ox|)�'�?hwL:�|]��"���Q���Q@dAS��r[C��dh���Aē:0b�a`�ܤ\ qH^���J뱱�S-n>|.lh��Ag|j�G�"�U�\���?�W�;�lȁ5::Z���tp�A����������^kT;��ٰG~Fd�����h$L��8QR��m�����6�������4�ӝ4��·�� 	ⵁ(wĲ����K���.�y�$�X)��7�Ϥ�/T�V�[lǔUB!�&Jr���ȝ�¬�O��AV�q^GX��GI��!�`�.!t����Tgྯ|S	3`�4"�g�C.�ݣh�ܮs����e#�vppО��8Y�P��'�ƆQ�S�-�(]8LT����,'K�8�� ��D�U�t����4��/KKK��Ի�^}�K)zk�\����`�dFV�� k5�[�Q�%':&��:�޽)f�<�'����$N����B+�31T<|�ӱR��\V�T�JQ�z.<�������A�SN�C���T�ţ�j�޻|
��gÃZ�ӳ��Ha��	�)c/P�)�������pd]�pJ��)#�"�w��,L��(CCC�V�,����K��|�ǟ�r�=l{1����"Y�cB�Aj���e�k�_( Ƚ )�~�:����C�f�=y��wq^�A�e��-G�4�,��ϖBxS�B���3���ݣ�( Ĝ�2ʻ�h*�2�����^�.{�8����GZ�d��ay���l8��Z�d�p"��'ct	�-Q5�,��x�KY��뾐�ݽ^��9|k�S_/��ɹ���{���$��2M���Cϼ���IRn�-H��0�	�yLp��K�L�L��G�썬{�)P��x�rؗF[�H�W���x�)���d	e������s�0|�� �4T�>*'�[ؠ|�%��8���C�4H�!�y$%%)ف���R���X���/��H�gr)�1��7�F��zZ'̟�Ӄʝ4�$�GI��S�{�8���P�A5d���b���=�p /5��]�4X*�	�q���06�DrGi��*�ء��ׯ�Lg��Ť�ro��"���utzv]��/ؔ��e�Z�,���cJ}}D0�B�V�8�"����HPH)H[�R{N�nv����!�/�$��:��Ũ�(�8
�w�=�����i*�ߴ�:�C�%a��X����Xʐ&�k.�3�p���˥ ���j�4:Ç��u��@en*��P"%�U�&��k�F0:f�MM1�s�oo��6٣^z�-[��X���KǄm��R���./�*�̅3 *$�R3��1����R����FV��8����sL~�u ����Xi-��&W��t�ƻ���G�+�$L���+0�2 �p6 �78Yr�� �z�=����L���R ����_l�q���i�$������f�V�ls�M�����e�65��V��x�Sp�˭���F���	�M�N�ك�����j-����޻�fw}gQ2/A��楋�%(إ�I��K����3cSRaF�GW�Z$�-_��C��Qi�'E��C��r�/dGp�ďg>�|P@��ۤ��N7����Y"�{��Ա����f6g-2]�=ъt�}��
�� %�G�(%*ߏNH|f�oV]G��I*o���M:��/~�����Y�~q�$6e�S���e[l��@�!`�u�)�-���$3����rV6��$����#C|&εte�ACS�ખ��o��EE�`�,�D���e���3�C�̨�r	�>���+6t!?����Pe�(I��xL���N �k�:нF7�G��*7֌�ÉY�q_�Z�Ih����ԝ����w�ܴ�j~�/��x����\�@�����KwK�!JTR�i��8#=����1���
U�
�JTQ�&�y9�j��s鄨�v ?�:�s#�8�؅��.��P4�O�k�R*�̨wU<\
J'8q��=���P�]���0�k@-O&e�m���Ă�e`t�gc�"����,\� �Ulf2e����۬u�	Ѽ	�|i��GP��ѭ[f��@��#���͐�fD'P.`�Xُ��U]{�_�<Z�2B:/���\K_ �������K�g̟�R�Q�^AH�+ʌ`����� ���ig�vcr!ː��k��Ƙ���{/B\4m�7<�	I�����;6�acc6ZѡO���Ղ��?<87��ǵ~�eûj�_�QM�!��t����9�3��*�jj�hf���_�X���
0L[�~WQ��1"�I �,��^$b}���֘dgJ��.j.�B�:��3�C�x��
�ٮ��{P�R@ca�a(���e~�O�U�Feˮ���\k����(���F��g�ք3�#e'BY�-:3�RQ-
>��E�&�0�,	8M�����É����GKBέ�_2�j��9���ќ��v����'���ɗ��?�e{/v������?��mw��d�jS�.�j \��nP�z�=��Ge$L�~rB���=���N9]�<�'L$S
χ��x���`�*�6q��q㘇>D����ߚj��Ṭ��t��a�iHJU�A�9q�s$�$Jߠ9���y�Ȓ9���ӧO�'�e:.��0��D�')�Q�e�-�r��v��O�y?L���`f��K�C��y������3�ǧ�c��q5���9F]��rxaNX�0Bf�:,�EB�w�){L��9d	c}W#����J�Ҍ���!�l�w�ЕN�g���eed��������Y���c�r72~�J�'-�F'�ݿI����L��c;� �|��}�h`7k>��3�`&Y�hӘ�	����!aPIn�����{��ѫ�W�l�1A�����BY,K͚��}��W�-�]g�xŮiZ�^I���]�q�dӀ�o��P�A�*=��Z�Q�wR�^��V�MM5��+��%�r nï4ra$B_�e�"W}OO��c(��k�Vc8���4Y�6F��V����:nC��r��a7�1	O�6!�\g�A$2����n����c}���]��!�0g���'6�!V����j��(pV����Q&��MV.�؍���k�O��	̏^��:
xe�u徥d���Q�ę����e�~V�񢉄3,j�M	:�:�QGU��G��z`'mC���sZ�W�hF(]�f���_M_�����l��b'�O�_��i+ִQ$ȔV���ӛf�E���Dv��*�f�iA�t��$l�����\r?Vo;i���pJZ��V�KQ�'���7��=���Z�Gܷ��Ct����w�4&nԩ�ET�۱�%ҁ4�ܿ%$"�2}�4#��3GT�A�n�5�[���}�1W@�˴.���T�ϓ4U����d�nɢ�$�����R�D��@���%wxc�r�ͪh�zAO�_?�>_ub����y>��2��$C��~p�|����xs��d�a����Aj��c3u�JRw��:H}�!�g�`�>�[;ѵAȑ�[��qr&&޸صp'׺|:x�~��V��}���
ebv(?�X�Pb���%4��ǝ�2��Ń2ԭ������N�RR����Hy�`��kz~�&!Y��$�:�B�j������q�=׊��BYy�����MuА�vn�48C��z4�O/���u�ܩ>�����Q����Dc�D�� P^LZ�3�����	��<��b����x��e�O�[GE�" 9i�)慺VF�w<�>�|�@���R�9j6|[HO8��d��ý��
�UZ�:L�+�?��j����('V��㇋ZG� Iyw�
N��/A}j�+l5�F��S ��yʶ���H~�P{P��b�͓1����FQ�� � ��m:O��lY`���F�ASѨ^�Fs� ?�s�3�Ŭ�-�K�%2=x�Z��}����L�g�G)�7��&���?f���}~��z~�<=�q�k-"G���p�.bP���|��q��t?�?���|@#CR���dЁ=�M����V�OE�@48���86��F���n *v4O{E�-$���bF�1%"�5+�b��GQQ�Z�P70��	��%�:?؄�a�0�H��\)�j)���^����F�������R+a!QQ��9jXw���dj�$�)�����̍��CV���6����Ys��Xu/�2F~��(�!U����B%b|�w3�?Q�y1T��C�
��	p�q��S��T�$x)Xdc���~�N�`��ɥ�e��ci#������Yr]��w�Г��e3#[,���0��ޖ����Z>~�Zo��j}�������/�fO�HB^Ԭ��|^
L#aN�H��˭"qQ"	�h��!���2
�|����G���q�[ެ��*�ܓ� �V�>�i��'����^~�'q�^I�[�dP�6��M=u� �xY�R;i�����iO��������!a���R4�tP��{f(@�rܷ����ruu�e��v�SG�K�xa;К�{�*��
S��;�^T�������z���T��3]F�x\R(.jqd�L������qϛ����#h�pT�X�l'���O��0q'�Tshη�7�t�愨�X�*"���/��89��̰���;o�:����1$�"�$o�R�o����؈���d�බ�5!,�>TyAi���Eϼ�t��W��~��<�؂+�AaE EMu0���]Va�/�M�
v܄\�f�G���b��iEMk�������ś��@�%�\������9@ǼQ�W�P�(j�DW�Qȩ��R"���Y�'�i�$�N���C��'8F&����O71���"���ۗӖ��!����s��Ejj�HϢ]g���/���J�r�[7P��Oqy�&�NܽZ��T��6m�Yo�5$	)]?,"][a?�U$U�J!x�F����T�8��ϑ���^i��lHp���
J�o&V*Ɋ���UӲ�&|�0�ϲRl<�R�g���$������^�~���O���c�H��nG��[b�Wm�A����|��k?z���u:$�j	^�X���!٦�+�� �$�Q��>͆/��܏���
���Zj~��$�Kc&�6�~D�7�+�5�g��U���t�2��E�wDa����v�sx����d^2�k}���"C|�w��o�X�.S{�'�O˝��o4�6!��w?�j���+}�����d�W!v����H�֬��ƍ����ˋb���|���@�,;�Ѐ���:����U ��˿{j��,�� 8����Y��k�i.�޹ÈK��5�:n�7;K��Jh��K�Be�ż��m��� �G9ͯ�y���牍�}~�k�ٱX誛��uCߒd����,EY�䔮����� gW�X�_�ς/��N���4#���4݆9���h444���M�X��~;���|��RE�44A?�i�=(��x�D���2�
���},Ր�$�uA�M��·��(�zŦֵ.qВ_\"�S�v�X�enf}��˩.���7H���|�_�F�1�98��N����X����2R����c�\���oݳk[�$z�!����S��v�`�P������fY�/S9�eF6�T��\�y�-���2ts{���o�0�צ}�r=QӠ7�x�f	0��c�M��E(]�dF�./�H}w�\:���e�����!99�Q���bw�����v	�j����<�`�X�]����Q7�p���_���\]���
g��ӈ�d�t�(}daOk��PdI l�0��bɂ�)XB(a=��b����K!X���5i��,�y������ٺ_I����p�Kߋ�'&�붺<oe=P<��=\�.�:�($h������9��_X�	V�����M���+����[�����A�9�T3w /�*)���5Ð�Y��օ�3,�G6xw�ɟʥ)9b�~7�7OD��Y>WTJr/�֗ΏmW2��Ď&l�4e԰j��f����p3%b��k����K��T�b8��-7s�0�h�l/F��сkY�0��@��Ě���	)!�6e;�ۣ�������#2=D�C����/do[;��/�����>_��=
>��N��i����C�I4�%�"^�m<���\��Y��Q��8��d�M�h��T�vSV�t�-S�L�:L$8�Q���ӓt�S x����ɤ�o��zd�:4U|	*Ҵ�z�z�O�88;���a��k��͵,(S�:��Q���)�����*P�j� >PFcَ����T����kxx/�9���<ߓ+T�^�8/_0�k<��@�؀�%��|3r��|��\;���X4E>�駠�J�H�ԋ�1��&;V׹~R��^xhh���E�X�Ҩu{{>� >��e��S�v(��2l/B�nS�m��៝*;�2����|�����8�0|FYVlԑ��ɝfؕc���G1K�=m>��L�ף��g��v�������	��DW�s1��(C�k���VQEvnH�b���Z�����w�9�������;�I��;;;�#i��eeI(7��yu�t���<�RP8?�W^rF���������������Ւg��8J�4<fbT�b�s�!�D/����V��J��@m���v�Rrƈ"�#���ʤBS��IмƼ���Ǿ�J�o&nO5W�3�l���3����f*�w����tD�N�<���(�I�ءs@R?2�O���;/�tb���A�<��C�X�T,��J�r�-��L��_��r��� /�Tr�\HO�p����/w�IO��8��]YP)�y�ʏ��r�A���'����0�h������j$�dd%O���hc&�@&Y����V���@bk>��sO���f1~Kb����³j#�5�@. ���������$�o"��G���.t�#�/|�:���셨3Td,�h�[�+�ލԒm6��Ш�,xp��%8�>�0��v���݋>����J��N��R:P�0%���\x�X�ج�-/�ej�ɨne���q\C�Q�Íp_��kA��s~�'B���J�0b�~ ��_�g���.=5~��F��#�#¥�k�=��#�p\@� ���i,�����X-j���{OY�NN7k��y(֌J��p\.�^���-ж&�@y� K�خ�ϻP�������5�T<?�V{냭-�A���KC�`�����=2��n��Y�Y)�Y���{���M>���e<�@�:�]�/�����7I�?/M/z��)w�����n&)���o��(ϗ�Ŀ4�p��ҥ�~�P"����L0�����L������c�K��ԏ0tt�]\�T��O�̔���~�T`�m�N�VK�^]t~?]�I�JP��|����;�L�}|q�k3�����ܷ������VTc�:c��_���>35B
^c%0�\����F��(��i]�n\Q�[nk�D˷����/��5]-�#��H����"�F|��O9媽+���SF�����#��}S�_�d��S������<Bꯢ��޲��5��>��^���8��6;XopO��Jhv������xل\�5hI�khb��D��`/�)J�3� ?�YjЪY�o�d�Z���q:�$Kb�������%��_QI�W�?�b��d� �g�<�Љ��'^�|������~�P	a2;,�� ��B�P������;��4��!���hS���|Jn���CΛL�U����(�R���#JE��gvG�����x���'�D�½C��B*ď%)+�O��O7¦ի屬��;j���G9�`��_:I���hX���]������H�of�0��u�k)��A;eg�G� ����������QH��?~���}�m��~9����O�#gg՝[?݊������=���K@�x�a�nd�B�h������"���Kn�k�3�_e����y�}�Y�!y�L�1���&F@�
����xկ=*�>��EgD�F;�k��ʐ�tV@�4S2p��ӯ�@��H<�A��3c�>�,<E��?A�-&"\ 4�A�L.;o}�[S�M�_�P5�G	z�=��3cEՐܺ&�B���c���o�x*�&����ȁ�l�mז�#2�a����U�SŪr Y���r#??���C�HK��ߋ�����)��l����:/]i����I�l�iÆ f3jyt��*):�S|�� >
sD5!>#%��V�!	������.,ݹ�	9y�Ū'jM�d[����66/��2��1�j`�P/EA	R�_�Q�ի��&�o��ƫE�ѿek�3޾W^����#���S5���v锔�8��.항�h��A��9L���X��7U��0$��)�:ɍ䬘���8�G����<<�>}���2-H��!�n�#'���Z�\9?e�I0���G=�������&�v������0;+�g�Y��s��$z��|�����r������B�u��9���[7�ǥܘ��|����oz��{p�B����BU�:��#WE�pY®8�1z�r�!4� ��W����n7��G<�%��o޼1w[@��5��v�����C��+ zd�+��3.(`2`����I0NU0�Fxu���Ʋ�u4O��|ʘ���") ����{����+�nm�i ���p�މ��hy��+�ȩ��Իn���p��K@O���^J��w�xӐ ;V�Wk?c<1#��{vr�W�o�vV���0�xWة%F�h|�5�cs�s�m� ?&k�&�,�?�"�����)�BzѢ����;����|�5x$�=��wm`�)cT�bS ܯ�'=���/gZUz�K5��}�������(=2{�IFT�^�f��+	�/�7y^Z���Ӧ;my"�7R����p�>�k����?�{�Tsʲ�X��kOb��d	�z����1L�Jv�X&5��ۥf���O=����~��x�.f�˯�s�f"� �:�A��mn?���E@AH�^fal��=!r?<��
��Q�Rc>Qr
��G�G�_��b:��<���/g�L�G��x5�'�ƥ��|��f�y�Nn��`��
��{�I�gp�C	0��3���T����_�WD�t�/������S�k�sn�=�%�0�X�,��{a��ҳv�8r�.b��z�)�܏Z�m!���g��6����Rw�:���!��MCC�d�i"g�vs��//��J�_@ܞ�1YNys�p�ܧ�����7<������P����������R��z���D^Dp3R��=���fƼ-R�d�C��Mc����ѪR��/����r�)l�HÅ'���KA_6O�^��M��섄WF�I)@��+ڨ�86�:
�Bf"$T�9&&	�t��j7`�m��#�yeyJbӞ]�j�=|�'���0�pd��^�OKs9ա}��v���^�\�V����U��bp���>;�~�x���Ґ/���Pn�?�p��YL�;k[#�s
�9l����k��+Z:Z�����a����B����!���=��K];˭�F�M������f�>�\�]��m�{��:��10!y?����x��e,�%�[�8&$ ��fT���U��8��L�k�t�M%�͓b���D��ɹ�&�[�U��t5�SS�-\�c,Ap�x`$�����1�<t��i��r�u��ЁA9�d?�}o�'{Y:*�B�)w�ػ�1�K���$�/?~����kC]l@�)F1��| '322����ߣÜŽ.Z��|2����a� �x��T����{O�!���4��D�=k�:��:JZ�u�Fx��Ϟ��ă\P{�0�%��:����T�}S����)���\���t��6���=�:��5+u�۴�|��=g�
?�6S�#�FC�H�`�зT�<*�93{�ѩ02�0�ʶ�C�Z䫑3�}s{(({�<�[m1����c�dL{��ދ�������r�Ĩ5vИu[��
��FF��&o�M����A�Hp�M�Q$���k���m�I��S2(�V3�uY��O�4�۽��v�L<���y��.j�|���@(�WYn�����(���s����P��EH���F�z���Pi���B��$�ǽ��S�`ڍYM�|2�]lLxhsw�ef��Q2l)�_��x)��c�\��ɾ.ln���(++��eQ �I�tNOW0��ۈ`�9�gn�%��AC�ɯy�yW�0��$�yh�.����SQ���ȝ���}�eϤN�ߍ�T9�K6Ӹ�*|Ã���n&k���8~���o��P�*}��b��;�HϿ']���k�n��_
T�R����@��o&a��I�����l	,���y���B��&_Xp�FK��ɥs�! ��L6|'U8�y���t��D��޲B*�jBO��%������<��!V�u���kZX7��L���R�l<� q�L����������qprJX���A����	�m�
ϻ��������4�^�P̮�t�KN��݂�/\�����V")�95�]Z���G�D5���&�hBΧ�o�>��$��c\ڕ��ڴ���d�"�A�S���{r�>8��3q�v����W{��
�����gy�c�����Ư��#&��#�����^�c��Mk�|Ng:�P��[h��P>e]r��7�(��f���&�]r?/Ny�v����+��zj��X�$Ӝ�#;7J��/�((�/wƇL�n�7���喤���
�$�O���y6UD|�=K�5C��P.d4�����$����#���.�����DInmz;���Tsv$��߿G���Fw��Z"�F�Lz�6���-�7#�y�L�?&�Xd�u7�5;�{�VG���(�'���pB��V�l���ߧ��<L�\޿�~�~]�Z��}�'�!A���i��Y�a08�F���.ȵf��Gh4���\qGom�
�Ң����e8�Eַ]z�M�{β���`J��˃�A�+~�z�|C/.�L�A��S�"r
+t��&D��]���1Q���d=�fQB�%�����h-O����΄z�,��TFa�y�#q�B���݂f���H��S����R~�苊2 aH�h�j���R�v��l�^����K-���?% �d�b�9��{�*���-���@�r"X�@�K�E4-5�?'��Ե��+�~#�tѭ��#�^c���=5�^ �K�|��p��i�w�%F����T���c�����%��YbN�+�����s������2F../��1�ii N� �#d:۵_Rh��#�,�-����c�*�́�7����X�������'q;Z鯝ƞ8w8�Q���/��<�XXa��F��ދ����\jr�0wf��Å\�n5d��Q�r�&�+���,�'ծ�6v�;�c�f��!����j�N)�~�:T��0�ڦ#�,�\��s�[�G�%&a`^�`�G��l*AY�G������Éo���[��9�?b^�|�\��$��� ����}�y}Vyۢ�0�	�r��ύ��?�Bo��Oΰ�)���p�L:�%�o2�����ͽ9�="ㄎyt�J)w	�Q
�V���TS�����!&�z�;�}�mm�8ߚD�c���7UXM�}3�b���55F�4��R�ڿ�<��I�?��b�T�_:/�[�d(��h� ������]5��e.d��>z�qݢ���>!A�ͨK]���s:@�� ]]EE��C6�o�:o�r�3�v�g�U	�&-�Bf������J�����V5����L�2_=ґ�W��H�g��?og:��˚��������h�x?�Z�D�#x8GA+x%��
�'@�.�g U�e��è�"*b��p�<|���8¤ ,�F"s�����F!*|Hf,�u�V��*|�0l/�P9NOQ�W9�b^$!�J�����7Qlff��5/�\̐��`�D8�J����̀�*�{�-Fl�K�Ϥ
���)³��;#&,�_�,VXd��k(Mbs�?��`���R�M�H�b�^��
�D�>�k��$SAn{=��) ̗ށVR6�� � �Ω4�:À� �h$ڊ��l�[L�]��?���`�󃲖cNmt^7�,��r��6u�R���h.��5r�u7��eOȂ�1d����l@��/_z4c��3aVOZT54D�uui����^&��QZZZQϗ΃���P��"��K�S��J��?@fe���Ȩ�#-��ԁ���Ϣn$�R�5i�A$G1%�q~W���Rb�y�Y���&��X
i]�?��1F`/L��g�{9��"�Eg=��l�kL-�+�Ǥ8k騊�E�wЇh���Y7V%�f��Vs	uu�;`m��-�`Ow�(�yS�~t�L���(�1���)]�f�ɿ&�j�V!Ҭ����^���n��_{��j���Ѷ�#h�7��!�$~�H5���7�7y�o�~}� Ht��.�{!�K9���w�fh�7� S��f�e[l��%��X���$��9������偅�kG˭���i'V�WW��@)�lx����J�1���"]������K4�q-E�bQ&��J[�ᇭi�;)�ͺ���ʴ&��|�9�R����ei�~�6� �$<U>������e�-� L4����B��H���X/��Ύ���@?&�s�^��J�Ga�6iV������{3�Q��h���Z����N�I[�uO��^�"�L:)��!����!x�q�j�b��+ Z�� ��O(�S���a�︦�<ۣY�L�\]�R�7���r4e�E.�6Ʋ��N�،,9�ah;�f�������d�(�B~lp}t�h�L�"cR�tF�W���=�~������B
=f�w�}
Q"�Fޔ?�t[rJI�! t.����O�e�G�����Z�g'pAd��Lz>Ap�jk�A����3��f!���&"(@�\���o��~������)��C���|�a
�kB�Է�1��$�����'�T�O�؟_q�-f���V��!��$���-�@(���3o�4g�CHM��f����S/�{Q~����Y�W��"2�#�l)-2����e"�ɣt���q��>��Z��.��.��W�\CIp���1�'Cq�C���PcE��������� �����m��oCz�Jg��貤`��pS�����	)��us�Ν��Ǎg*@���qO�<wg���$aO��&�=�wJ�+�
�Pz|�nɦ،Ua @�[2T9Kt��4��ɇ��N��B��$	�pp��F�|�8��MJ�j2�r=�W��{|��ԁ�����|�"�tlLA~@R���S�߿� (�yCN<`j�/_ ���̩}G�
�W�k>S�{�@�&���fH�τߞ#n�#��L��!���U��u�4A�a��o�h7�3�1������m�U;ڂ3(��YX�� 0�L�5�a���O���DD�R���k��R	��?�1:�F>MhMĹ�dX�n�'s�����Y�aD�`M��$Z&�F�3�2���C ��7S����3�4S`��׻?�Gz��x�t�C�s�fc#hN���p�V��P�P]Q�6}>�Se�)�0q��\��逞�*��e�+|PZ�[�`)!�j�I���⛸m=~��#�B�|/67��~�a��!��G&@�	u�5�H�i�J�?�%RS�f*�/�;;������E��<id!�{��$=gj)Ĭ�(Y�y��%TB�zZb>%�-��d�3$�L��r��V����P����!S�L����n��i��s�����ZƞU���@����Xٿ��Ǉ��[M��\m�gg|��a"�$P�^!(h\�����o��ה����~r����@�G �-��C����F��5�����"�DL�\3W[�a���-��	����DߓI0'U���~��Iq��/������n��/�����gg����^� ��ݐ���?Y������~�59��<ʢ^�����w1��X��F:9'��-�0��Bz�F�*(wGH	.��a�;)>v)赇`�C���R-Y]�����v����j��l�z�߽�~|�Ǵ�OL���!��V�Ғ-�aln]�Vv��[�O�;�TK�d0��}� T�.�1���v�ѷ_���~�T�#�l�t0�g�>Z�$�qG�穁n��{�Z[� �<0Ʒb��������s�dI��<H�;�}��k8K��w������e/B[�)�ɶ��cdbw®�<���]%��O3��gt&����P��NR�Տ���7ֱR������/g�;�`<���+��#�:q�	��t��'�ܲ6��E;�C_�.�3��T�AIz�r�
�*?iR�~����m����@��YB�
o�v�j}jLU8�{�ٽȫ�J�~�3%��8���_����Ϋ���T8��Ň�xQ�aph|"�	����Ej�2��A�'�,�	5�����(�u1�ߺ�+���HѨ�͏�����n~]��ˠ��Bo���3�,<�h�{x>�k�g���M�����\�~�zQ:���),�Z�.}ǜ�m�6����"��Sʺ�n��2󋭭N
u�&$1���n\~�$<�ΉL̗��+��ՠ{�&��`j�ʅ�1��D^ѿ.m��y�%[P�5cx�*�J����t�d��/������1���=����\����ܚ����H�(��*���mD���W��2�7y!��KZ���f�So�'+\Q�~�ԝ7�����:���f���2[�RI`��LE�>D����h�b<K̠��v9�G�ɤ�ȑ!�qO���<f�(.���{�B��X㏵�h�1k�c�Iar���޼��´��v�5�AHcI�ѝ甎;�<�h����5:�� zoPAz陹O`��*l�R%��<R�R��Ϧ<��*qy�5��A��v���[һ��9Η�p>���`>ט��$Xp�<�ry��p3r.}�QR�	HP)��̛�S��t[��jm�A*�d����]-Xa���4�e�RV�eb���v���_�4i��KN�њ��>A{#�"�h���5T�wwFd�H�!����4ǐ�0d��F�&��!<����/1n�^���WdI���Rj5r��L,¶1B�1BpՇt�~�MX^_�c��&�����` i'��>��=`[/����R��@��Io�^�t>��RG��)T���y)7����؈/��Ã���&�o�M[����^�q7�ZD9]*���=���꽒�����u�Ag4��Ih�<��m��K�[S�����Ű0�������!�:��$���u�B�1n�2�6uT����eÍ�8k��0�<�|�Y�ν����ge���`�P�Q��t��u{�����,��j�6�kpw-
4@�ww��P�H)��.^��
šH��P�hq��޵>V~&�̜��}�g�L�3�#Y��GC��v�8���n�4�L�k[g���I��g��'�ƃ�kf��� ��-�[��+J���'�5�]v��P]���`x�0c�r��P����퓉`��S�����c�eUU����[�-�\��yI	�q���=��~�3CC�F��,�&�֏�� ��H
B	#�6EDD���C�!������b����w��]���gM+��7?>�HJ+�[Xv?=���u5$�A�S�����sR
4hW�6��\=�***nDn�741��\�Iiյ���%�q�xmޓ�V.�E��?�����.�πq�9DK|��Ąӭdf)�B���y��ߪ�EH�q���.�<-��a�?�^ֱQ$�a�<t�2�u�Ƕ�v?n�
����M�n����6����Y��Q��ؖs��ʶ&������O�\���{��7Z�쁔J�:ۊ~o��E��SH� )*�:�e��X��?���c��C��See����vD��y��`��{��L�<��I���R��L� �4�����0�.��\$:���gY����������r=F|�[�H��r<]���qRbPپ�>V/|a�EE�8���OL_����)��a��g$ƞ����n�H��0}bD?8	*/m׺�Ɏb-qS�2a���}3�0���q����R�H����jȋ�4�D���S"g���{{;#��Nj�u�Cg��}ࣣtu3ds�4rG�H��!�<�c:E+���)6W�]_���7;��u �1l�=&?����g��2U��S��uV���c��t� 8}���#6ö �#mⱝb�[q��nsALo"Mv��k�=���j��P�M��!�\j�佲R�������Z$o��wy�JH�P��5�0�{����7�Cs������0�;����7�ɖ�gde��M!����#<�Ud���ﰻLKOW�H?^y���B�rL/��j����#$���e���A�܍��q��'����`!!,)5�9�";�:85�S��F���@a���?фR��8����٥t��:������#�F����zS1}�t�i���>2`S(�xʆ���.���x�SM�K�=�>>�\�'�uh��m`�uV��y��}}�:?t&0����!uQ����K��^]�*��>�C�%*�NQe�,\<s㭊"#�B2��U�E�&��p�K BV�g��㇗KÍ�G��y�c����-���W+�Eh�j0�`jh�t3�i��?bkȌ!��t��n(Ε9�|�gy�1���b��J�y�M����%P�׮ޚp����	�vZhG�����b�^�WG�Җ�Di֦1��B�|c�rs�3I�2h~H4�{3�ݞX�5:�/�HQE�(i����l񯑝��a��'�n�h�
g�x&C$x��K����?0�o�Pk����I�ƾ���{èa���� Nc���%nϳT��#��^��.L.ab'���	�7Q��)�a��$�ORX�o����~�j���E���7u2���BK��r�����f֬X&����r��;a��Kw9���1Y��!�fN�hMb�c���?v�T�����P+��nʍ���\��@�����z��<��l�n�OT6���e�nv�'}�`�n�W�-,MC���T��8Ҁ!*��Q����pP��q*����9s*��#��/NV}�r�v�f�`��&UbD`�-��6�z���"7�����UB�
ql+kkNcf4��� ���9��e8M�
����OuM]]	��#5�� ��0���/��8����L�"h�Cf�쩸��t
��?��j��>z{[̗���ƒ�!*�Ll�R��Xò�3��p+1�1�\�:���u���Ks�0:?���0��c���\���{6��M�V%W�>QԶO_�t�t�J!1*4'o�Ɠ-�M�`{^Lnr)������kD�c>�'��=�ʑ��iMȆ��DY��u�#���#��Z�/HsvD����olg����?�hV�������\bg��5`?���ߌ����g_m`�������7�$P'��_w��k�ڕ,^ Hk�>aݒ}�)W6�T���9�ƦX +Lp��q��a	deeU�`�0�j��W�Ċ�ź�D���F4������ YJ�]13�����@�ש1���a�T�q�ّ?��6GK�􃗚V�E��v�WOo98�fT� `N���=�|l�p͇c^��fe3G?j�a1Y��H����CեMp��r1Ŵ�W� ���@Izx����RN���0p�{{	0½������hƗP�}
䓐�
�r*�NNLlw?�������=!J�շ�E|��M����kw�Ά���w`�e��ݰ�����у��i�R�<���R_���=��6��_����r����u����8�̄��c_/siI�R��/��m1c�&Y6/��(,��\�]`�d��@u�)��Х� W��:�2u��و��X�)YJ,�� ���1}��z�^G{���v�O�5�M����T�.�$��5����D Ɛ��-9��߃����g/�>�c���<U��(RZ��E��^�;���k�e�(I��f3+b��&'H6s���rqR�]��@J0�O�,,��5:�J��u��Y.m�FH���5��Z�cM[j��O���;<��6�.��qp��Vz>0��Ԉ�_
�a�ྍ��|�T�x~a�K�sG۝$P�C�I�p� \���A���\,I_�s���m���
_,����z��<B�����P�[��nA �9k�1exaY;E�P�S�"�ǿ�v�t��9��A�З����r�>x���쀨�.�eȒ�m����d�a�-)=�qF��;���/���	!����>tv*�:a��������w6��V�/��%�9��N�?_����+K�t�H!� hZGN\x�:��7�҇F8��Q��Ę��5��7��͇�a����z�H������S�RLK����|�G��L]}}��-�����3ܹ���~=��EJ���kx
�i�A�E��jf����M�6��
�������2���<����nn,�	�Q�n�*
�N����}�%��ɼ�ɉ|�c�%{���Np���Ք�~���=J[����ߨh�v�))1���2��p��U5E���٣=�-�B<�F�e\]{fly�%�h߄��X	p���=N�ϸ��S����aj�������������f�-yʰX��qPBݨN#���t���$�ʂ�o=x�9Qy/�@�?�K7A*BdH�� z��7t�{[t�oOc��c�L�m�\3#3S�D�(]������7Qg��1��Wk�����y�wd�bqy��HC��� ��w0p}���a���v�Е|a$о�
J�mL	D�Y1_5��?gB)C����ց�})q<uѧz��\��߮��KC�����^�8F��ρH6��ŵe�2뤽/�5�{T�����b������2+~��㿳�3`��������E b���A��ww|ll��q�NB�@�}����B�o��q��^]���eؤ:�D�,^�:��SƝBʞ@���TZp%�qzeT�Xi*�k�cH�ڕ�,�%���p�i�&a>��*W�P�jcނ�� �����ҴГ|<A\����M	�V�%#7���
bǳ��j�M"�-��LK����B}kk�gL��v�=��Nm�@��c�	R?!��^�'��M{�Y�m�K���a��L�������,'� |���ż�4�lB3�2����Uҍ�h,�PՒ�p�П+3������8�6$��C��6 ��yF󥥥��]����"G�+��MCJ쾂lXU���.��B�@}6��YƇ#G�ZV�ʦ��@b�/��#t�լ�xӇGj��+`>��uW+<�l����t)�v��`$�k��gk�I�#۫��N��n.�B���#I����K5��ҟ���CnГ?�<��|Z��W5������v� fм���l����������e���_����#�UH�����E] ���;�����0��9��X��y���~Xl�p:�}��1242+,�h�D$j����3�'��;�[&�0�v�>�ܵ��褂>����|�q��u�L%����!=u�M4��EI$@�9�F���0��*�]����� r��SII���O���͠~�X�0o"� �7!��8���DҦ��'���,('���3����I��Ѯ�tC��B#t�D9-��MF��3�6����ge�����Ί�]���l����)~I<� Hz�'A1r��oi�����g�v؝`�
�++����<U55�-�\zr�?�4�B͋ J�vf[����̪�fRj���7�c逕��������2B2�c��\x/!�NĠb�м�f%O�_�������]뷾@�@��c��?�_ V�>����m�����d)�����@���
#���%.3��O��o����@����*��ۃA�*/W�@�� �Z(ʞ����f-`4bjD ��O�Z
q��m��&��B���V/'���������b��o{��u}�j�MGE�ȕ���r�b^,Z�,[<�\��i{3`�;J�9��kOѕ	Vm�p�%Ո������(��	�y%H!Xi	[eC	��D�cu#����������_�p^v*�
ٳYR��"�P��R,�w>e�tt��Okj����Q�;K���:`�٥b8���7-�Aq�%�G�y���C�+cݸ�pc�(>~L���U)���c5w��Ub�i��sdDX�8K��A�Q�<o��6�,<����^׃$áz�v���E�֚"�P<N
��V�s�'5�֠P"����WSM[q ;`Ɯ���i���S�\ �Z\�`��A�	���Ңj�j�J��q_}���xX9V�qs�H[��x;�}�+w�����9�)-"�d���̧i������֘���xJ�7�(����-�5����ljFR\V�nJ�X�+@���^�(FJ�i��H�%�-���<�Ɗ�d[�r��=����}���9�N�������e����뽿��S�^�#S�J��Ǭ
��7@�j�����̾(D����T"2�ԭ�,-�Yx�[3���V�!�<n����nh5�	��Ԙ�����j5�("56��A[HC����]J�� D�?D��'����r;�q�?|s	%����ɈmBd =^�L��`�x �F�����P�0�o��--ҵ4�s7C�_�*֢*]FJ�iW��#h���WW�o*pWt�j�ͼ�	#?*��η*���f"gW�T�����*���Ŏa[� Ӭ/%���%W���@�ŖX�ِ^u��=�쉨ѕ_����7Tu������0^�BC##��HIP�yѴ���Q�S7B?�ԝ�E���RO�R�,J��Ԉ���/��ƃ�wA�h�D�
`&�4Yc���>1��2 !]$� ��Xx����ѥ%�wM�eCY���-iG,�T��F�,�Rj��^��?"�)E�i Z��	�~ZQ��4�Iw�a4=d%�4�����/�.��aA�z�j��}3h.M�H?�w��N�Y;�5bp��!zNc��g�������~��*߫&Z�9�����S�¸~݊-�?��NW�N�N���Q�v7쨊BC
Q����ܷU<�^H���~�DW���s�X+�9}���eT ��z����[g��x�*&UCa�7_%�GݗV*��$pq�����k�y�q\7;R��_�mI�Ч���94���V]�ҷq?��dm-��%��{ �T��۾"i-��\-ӌ�_sZ# �5fB�evF:����^S&n��ܗ��ӲI�]�H�)� ��4� �f�+#=�(�t����0����pߎqُ����/���-*������4$����qM�r���}\���b�����ӳ`������cZ��X�1j;��N�=�?qz��HB$�q�8y��0܋��g�h�-%r�k�j !��SK�pҀ�VȪ�>i���n���}׿�s�(3dKg
����+r�P᪋�K�:�t���KB�lhG�jm�|a��E`⵾���T��A_k2���s�$}B�;�NF
�u��ͳBg�^�&
DKb<F��v�և���X��m��������m�f��s�6,d�"�%�y�4�u:��Ⲿ�����,]�t�� ʢA�&+���?��Sщ.}��݈{.�с�Ç�fM���Ԗ���rI6{�g\J�P�����2�866ӝ]V�]SR�;j�C��xIh�����O��É�Y䏮��ȱ^9�YL����}��O4���P����G�)��ZG���*K��э���9�h�����J�Y���n�kۋ:�$67lQ<g:d����sگ��5�bZ�W�e���Ю-�����}����@"^��B�uɖ x��|��$或�cz���_8���[hAf~��x?�(��JU��c~Y&�#g-<n%$1��K\$�bln<!��i[I��ɇ6��1p�3�ES2�`�M� �t��W�ˢ����B�5���l��_���X�B�ʹ�׸�o�v$%~�؟����:_�C$�L��R�-��xښ�%��X��Ķ"ݵ��u^#տ	�ݹ��_�WUq��*�3��\њ���J6S,����Y�������#e�#%�\>�Z�H��*�}��Z^!/�B&�7c��Tp�L��)Xr�z�lZ[D�i�CV��<pr(dǪ�.M�h<h�UQ!�}s�"#�Q��;�n�N�1u���np�.����TM�A(չ���;.� �(I����$�@X1Dռ1��`@��TJ�t�x��S��)� �2&��������`���������!W����N�Q��"�����9�wo�@&�H�f[���S� �`��4ܐ���b����^�!T�x?y�?2�@�'zSNz+_���R~&����9bx�l����<%&k����Y���ҙ�x�ѹϵ3��+	����d�Xq��Td�Gj�W"�9o�螊����� l23���_	V�V�ލ��}}�p6L���of X�>�n�S? ��*���b��74�e�շtD�1Ş��~	:)Q�����4����5r��ꥥf�)c,H�������Ͼ2p�z���W��VJ޷� 2�Ya�C�?e�_S6fE���IT_ƎXS7�o�Uk+|�'�ؔ&�T?A�*s���b�5�	��(�`#;��z�'1�`0j��IUOD�MJh�dYe�!b��A��i��U,�&�$�)ȥ�b~�ٷS�eI|D���<r2t{e���B��l�O��m��~4m�^Y�c$U�̶�;Rw�Ҙ�/�k-l�a�k:R�>59ĿBY3-����DK���ޔ�(~���r'�*Sg.��|f�.n� #�%"2��%�</n`�
�bc�#]P�L�F!��'}(߽<������ً]Qb�J���M?��~�KE���Q�oj��)z~�#]�\��E��`�bZ�o��f���1G���+����]&������?��+���6;�df�v���+X9�ϛ,�9�O���6!΀mH��G�`�gE��	�Q�<ЈCo"����,�'C��#ii�;V���Oկ`IA-�+xloC��ܑB�qzI�� �F�K!�F���M��y�t$b4e%�c־]�l���-S�8���Qk��N@$L���NJ�q�䣗T���E�V��f[GQ�Zv69r c���ݗ�Z~����[���T�$@�w?���q�Җ�r�T0O	Z]5�d�.c���bLg�.y�Beb��̂+R�c���FZ�d�s�(L���� ��Ȩ7�"+��5�Կ�L��"�i�d�2]"F�S�A\/5�/�쩧�,��d^�^������T��5C�%�`z�3�`�^ݓdё����VV��3(NCUϭܛ���O1�����'�J#����ֻ������� "���'��#�Ddt��R'��w��	�)�j�ev6��Q�`C`��c�hǸ���ˣ�YC$ųbw�b����R�,_�:9�tԘ��v]W{�dOn.7W���3O/$�2�ے��#�:@�|�L��R%�f
��P�ϲ���Z���T�C=���T�t�4���<������̯B�m��	�%!Xt�Y�L�Z00)V���)�N�\�}��76��]�
R��/��#����Z5�a�dD��S��<�s�W����+��:4�s��\CU$8�<���r֑�HP�9_�E�<��wQY�ӇXꡠ�2�I���G$8_���My�|6�@����,���.B	QO���O�ُ�Z�3�
b``p�}���g�������96n�6}R�bm�j�%3�K��x�"�f�^;������%"4�������������`kаY[J0U
I�Ӆz��+*̾�=�\��c!^�X6'�or�K|r�HUr�V�d*�aH��K��J0,פ������I���ї����_�(H��7���$;��}��\�?�CXW^�#��l4�]?��lV*�O4v-{�v@���bM.�1DO�uΐ��
� ��&��~�]���$�MzmI}����A3uw7����D��Wo���&�Q:�����mc������g��U@*s��Px�5�N�@�y������X3��hE��f-�g���JK3F��DX8�&%i'��W��3�%���z�{����ե��I?���`�}.e�S?��T��,\���rSoW�6�r[���3�)VG	����02UJ�pB�9}-�m��aܺ��Su�N����a�P>"��#{��H����Yq�d1����h�t;����/�X%}!�c1D<�A�?σ}�q�����n�o�<�ꇝw��~@�r<�#t=����70Mr ���K���I}30�!�s��i� Z=-���Cc7��a��=����r�����Z)��6�Y6�C��>*Q�r��9G*l��\fd�'ɑN�7�B5��p���]Az�XĖth��Q��|�����}�30�i$I�4��b�a�da ���_�����f=�#������6�ʚ���Ͱ�oW���� �u�z ��m���Y	�)���h�ƭ�����s9"�X:Ād:P�w��k&��ه��%~Qb����6!W�fR�.�DJ&�P_�=�{5�8<-�?�R{qB��������\ޫ|�kt�0`�v���{UD��m�D��#���>|��[#�R��ʂWWP���Gϳ�pfK�4��e����g��<ޤ(X�U��Yo�������9'R7�J�ԉ�c�|q��,�[�4�e�,���9V���������p5qfHBX'Z ^��/F�S�β�w��)�=�_T�2�ԞiM����8ԯ�s�-*M��pҲ��O������{�I�qv�UGs˼,,S� ;�^<[��&�y��7yl61?�c$����e1����8-a�N�$1��Y o-�H1��wS5z�!
�KȊ�o������ E��\0����a���*��k����� 3�s�O�g�F����]:�1[�Q�ɺ�{��qI/UOiLTCˍsll�ue��K0'�v ar�S�3�����7����Nb�jO%�����v�q�l�.�S;�\RYY�gn�����l���Z��;N��)�KĠ���(�&��|��ڙd���T?VШ��P�����Lr��h������nC���;��)��]$�3���&�B����#\O�[��4���e��7�_��)���JhH7�GTP:�m�I�Ҟݜۄ���҈\!"U���k�l��������c\9�-Ɗ���q�Y�=f [9�M ���U��́s����@:�ߖ���MÜ��k�Fk7H��I�{��=��E�z0}dB�dҾ�?M���}��i3X��.n�z��y���*\+7 �A����n͇[|w�w:#�6@@�q���Ψ'�h&�ET�E?��Eݱ�K9;�����F��u�5�Q���_?#�)":]�p�bb�P	��{dJ=(ƊG�(ץ�ZȰe�{���ՙ���L`���(�����=2ǥ�ecʨAy���N�.E�%����Ƚܷ��/oY2�w�QUԅ�0-mm�~��s<m��D��IW�����=��ih�J=CCCSB�>~zi�?,T��a�db+\�zb]Ӹ�S��tY���}[+04Z�s�hs��ȯ���o�ӆl�<3��X�kw�J�0�I2�����]��~���C�Vz�i��*�;�˦EKc�}�H�Z�:�B�)9#�D���"	���[��Q*B�O��2�$�*,4�}Ng��j�M��O�,a�x��7��[���1�.ث��H�l��\��}"Ca�YE��@��.j���JiSUl>��S��qLn8Y�_V��?]tw~�������M���nu�:�A�T���ʮ����w��{��.$6��_�tc�o�b�jP|u�ppNY/�I���
��	+�
oKkk�\���zU�t����~@�~v8EB�y׶r\8m'��O�t�ޜi�\kLb�������!�v�?��=�����0��"��T.�`����!6�y}��FH5���}i8�hG\ɊAH���L8����iԤ����x@9	��sy6p��4�E��Rؐ�Ϊf�1��M���8m��@��p̦���I�(��,Ͳ�ƥ|�%WPU��?�I��k��|�S�:x��= #�;9�w|
�������>�s` -�0�n|�"��������n�|��I{d�ŨR����D���.4���E�:f*�8y�SL}��`�+Z��ߔ��M�H4���|X ����0밦����PҘrl����{�����돕fHU.5h��nlnޮ�����\��a��Y����,����� �m�e{S͋��s���C��cYf�Kí�i���){᷎���ĸ��V�]Bi��N�4�*���� +$�Z�f�ϯ�%��Fh����m��]���W4y4��	÷#�)*)��������?���q�277'}�)t��Oޯc�j�
�����
�w7|�h�Jb�3>�$�(kA�nn�R Y��k
��L�w����	=�A�]�-���w��~3�mn 2����,Eo&/�
\>�4������GBOh�vF����T9'�,	�v�r�B_e���y��S�nZ����'�U ��9o�����zx��G���N���&H�Ո�74�i�JO�)򓩷{<�����c�����ò ���6J�_x�7*�7N��V��}O�RVd��C�Y;wy��}�7����_�b��w��˒ҟ�n�{�����.Sr����ss~ׇB|J;��d�Dµ�E,%{c���@J��\��qP�Y_�kdp�)5UXS��񐻅:����X���k��Ͼ$��5��No�V(E�@N�+mΛ�/���N/7N�\�GT�n�2�Cr�-�6?9CCʣNp8NOP<74�>�y�d8D��U�����)3��KO]�,��J�l�ݸ_L����e^ǈx��5���8A^���~Hx�y*�6���n�㊂J.���ژ�5XR'��w�i��?����3���50�Q�W��RRJ�1�Q��sX_�ʹ���#���D=A�4��=[�$}��z;;.���gp.M�����9�##>��&�I���Im��5+�Tss��?oD�g¡h�i��/JP�������n�����:;R�l��Y�ڐ$::�U8��Q��G6��0�<h �x�6�_S�]�A���P��8����9v�����H�����r�Vo�!��5tn��nk�� X��W�q'�X�ڈ��e�=�mKd���k?����E���Ą��i0̟����:���Wo�۴��\�^ߤ��"��h�����@ܿ}�{��±��y=^�Ɨ��f��ۼ�Eg6J���%Cl��*w�n�l���i����<�2�=������4җ|�.?'N��x$|����yo����&zE���G��Ҙ��r�V�X/�o�Nh� 	���|-=��Ȉ=�a峏��^"j�f�E����{������Gف�颶�OT�>ء��ﻮ�|u���FyX|\?C��n˯��X�9�5����=����JT����ۂ2s )a*��g�<����%}	9v���F?���8�}���]��1�����OCV�N��*}]���V%��~����MK�7��]_vP�&A)��GK�7A4�Y��;\�:(��������ʻ@���ĊR%��4�+D�Gg�+́�Ҥ�h�ϟ�C.;Vk0��MBf��d	���%��F?i�枠��m�����]���|�拇����
��ak�	����FiWE�	3�"�i�t�c��Z���T+��orosQ3�7)�E�������:U�oUL�������o���Fd�!���Ꮾ.�R�J;��OO߮�u�iL?}�ONNv�H(�ǟC�r7B#�w�����垄��s¥������r�^���0(�֯����}U��?\�����8��/�I�Ӗ �Vԏ��2;��Y����v�Qvd��k�w	F�"�K}����9���շg���hŘ��[�ݾ�$h�&�V���oL�w��� ��̀A��VБ��6R����
j;�M�Y�yw#����ۄ��ܔr�Lh�T��g�W�-�w�枷�/T����}6�\NQ��I�A?$����:WqT�S�ZB%���C������<�A�6$�Fur����9�K �	S:������J���l?��­���͟?��Q@�)z=�	v5I�!!9��t�=ni܁�>)�E�M�d��A���y�k�wo	`2_}G��-b���P���Ӛ:ߕ�`�ڂx��Nd�
�p�a�N�1�=ϷL����x��8�.N��(�����F�2��f�E�^B[�W��㓓觊+���<���)^�D�i����̦�J������"��CC�O�;����׍O`,W�F
���M�;������7��4��M^�Tf��C�����S�����lɷ�׆��l������!�!
",<��͡��"�`�!g �*�#�1�F벅+��[B�v]Q�;�p�$|�����{�.�G�O��Vla�?X�X�;�g ���*	
���<Fd0�Ic�Xav�J�[�I���ecY4�'0"/�T:��z��p�AQ�u4�z�����qM�|̲�������Q]�Y�������/;F�Em��l�F��r���Z���$!��F�� �O�a;}�?LzK���V�e���лO���k.+��,t;k����f�a;�(Q}r�Ŝ�6d�AP*�_*���bɵ�����ٯ��E��ؐg��UG�M�"5�d���h��F`ƀ[��nzo�IO<�E u�뷽:1kc-3q�3e���3ݱqTe2�ˇw}U5�[}�
�Ϸy��W5���w���o<u�5�����0�1A*E��-��?��h������~o����P���Q��6���3Z��ha��G)�,����s%� ��h�_2M�s�s��G���H׳?�&���|%jN!*~;rv�4��������53ZRJ^A��9�av�٢��P���Ӫ����ɍ�E������.E]CB��Nvo�B���j���^��~��V?�U�B�����;_�[�j���w3cm�}\����4F������9��o��qس_������}Hz+���8�����~���翤�"�O	/�_���sj]��%�-�@CK����kk��B�~t3"100`NK�D>pC�&k�e��o�R��_�����C20X�\�LJ���账�ZZ��]��' ��#݇�9��}}��t��l���B&���B>��D!�m/M��)�3Na��6���ܼ�7�׌tݨd!v4Q�b�t��\�rf�!-��rcV�ʄ.��>�
&_��Zu��}�C�EP�6�y��+'�$�<���Bё?2� P�xck�y�9���?������/���a5��r#��2��
��C��{ޘ��߳Wl�|-��ho�;Pn��Zj-���ji!�Q��5�∉*Y�Sc�Q~����n����@��h�dv����o oP��H�ǘ*�Ԁ��R{��������<��ej}#����p���/��'	U�����$�'�i`�S��o�H�������5�����]����T�f�/GzZS�Cp@�f��V�0���]��ݷ�ć���6 =����xy�;ߊ~�{Z�}�R~y|F	��xW9��p֘��f�"]�PT���EU�0�Q�u6W0y��ސ	:l&'�M�oo���Vh�ߢA��a�����k~������w�J��Z�7y�H-n4\i]�5�;��C�^��)��:́���i�d���;�~�R������f��*��H��[���M��<N�H�hr��f�M�x�h�^��z`�'�;�$��g����Xu��r;�4�-S��q�!�<m���^�$�̄�~��鉸��3���S֌����W��=�7��K�����JL[c_��Ø:��м��ҁ�A�����'i�Ċ�{�����E���`�55VBMgǁw��E�,C�h����PB����o5�m�B+��+~����RE���W�����v)�<LMJ�!�v-�o%�=1vߵ�����j�m��_���?����x�̕빅C2�(_��ݽ1O2tj�ZJ�l���g���K��H��8��n������T��>�е�w�E1O-D\^�
��.XpIi����H����
#�lw�c��-X��;��۩�H�u�Ҁ'�k3P C�2�ĸ9Hb2��m�ʢ��%�#��cɛ�J�!���B� �Ző�8Z�e�s.�y��\Z�R����S�3��^�܌q��qƋU�1Ƕ{s+j�)7��6zm���œ&��#�T%O�X]�Y𵋺�!�*x����r֡_�_��8�T��y�!��j���������H9;2���U�}�����&6a.=���P'�vI�>;�c����J�@�9���*��go}eA�_����$2��!��Hqmj�a-�C��GWF,�U��^�BM�E�*O*h����H�Q�jY� [���Z�?�� u
���7����L_2�z+_�a3KA�_�-�i��~+������Tcl$=y9��ޖ;Ң`N�k��SB�d�cGm���ޖ���-��c�?�>�8�����3��m:�b�
ڇ�	XKV����0�^Q;��;���ٞ�#�z?��,.O1�FbL�&�)���J~�]�_\̰�<=>���P6�7�,�kD��}�Mܽ)'�+;�\��Y@�Y����D��'$�'�Ѐ�E�uNX]�ۍ�g����ŕ)�f�z��R���\@�PW�>�x�:�#k@`s%��>�~��{ݸq�,���uB�	1�[W�ʣ��,��UT�����i ���$���.�(�3
���)�]{��޿CWڐׇ-|��q�x����y����J`h�[������>ehݖX�s"z��L��bzJG.��M'�Ƹ��ݾ��=G�)��>��-���.� :i��֛k�� ���H�v��"��zOЪ�-Oh���Ɨ5v���U������o��O]�:��)�m,�
�O􂱮(+*Az(�pzi�
Q̿m�䍧����x'B/I�gYʲ����
��%YS�w6�ӽɓ�Y�$�P9?iA�---ӧ���,�������\̑5�����8���lϚ���TYl�?��w -���|�NX��0_o�����#Ȅ���#vtt����g�������z.��"���%ݲU-]��\��:4y�����=+�>�����x�_��н㪘c%0��
I�$��$(����7����݆����Ej��[?�}|�ᚙ�}�`�E��mӤ�c�Z��_�$ʓ[Kms1n�ޓ��F�G�+n��A.m3�p��:�oH���������CppT��� YY�_� EgMŠ�M���K�E�37wr�R|�Lb2>>��b����KhS�7��%�Q��떍y��sԗI��S/j��~~�'��c���]�D���F�Gn�/��lTQ��a}��T%��c�3x	p5{AWh]{U~�3�536��`��@�A����0eQ��7d�-���G_�@��[��v�Y��Lt�*/DX�z��|0�$1��a�#�w�S��&��L�_t���MA=��H���e�$���ܽ�83Tiځ�zU�D%�c�8�)��m���	&u���%1�b�?`㽑�\��?��>����`l=R��|e>¼� ,<�)�1C��K�.FJ����������O�"�p(E���i�-\|�O�D������|ht#$���nQ^��iǸpOH*j��핛����&�<�BJ��Ȉ�����D��VT�]��%O��l=�|�똇�I�(����T�n�`H��MX�h8�U��4�|��� ��P*�������#��������4R�VV�ͦ��"S�}>Lx�.m���,Z�L�/8�bv�|��<�h�ZF!#ƶ#
��!��$�d	a���,��Q#
C7��e�k_�*.\82 w�ŷ�P.9���q�W�2�s�N���<�W簢��@q8�����"ީS�����oj:�>���5�IH�̲l��>d�A��#	}�.a����C����z �)�<��5����d���2x�#1��s��T&�H$�4��f�pVV�Y�O��;��O����q��7MS`߂�?o�
�EE �햹�{�f�a_����[y�kJ���zYf|�[�6FM�� <��qˢ���x<~W� a���?� xA�E�$�kqcI@@0��8bط����fq�J|.}�c���hT���,S�\�u�H��:�~���	�J"�뺈��4��@��ak��}��[�U��V���=���:z����D�U�jo�t��
��4�H���=B��`�0h��(��VTE= v�ӫ�i�� ��	(�������"�vH^W�!�cò��蕇�V��KQ�(��v�!BX�'����"5� �X\��GOL|咬��Q|3������]D��t�VدW����ׄ��İ�!�DTYB���k�0�� l�N��6���,e�@��UN��*"�L"��R��Ib2GA@����)�������A�F`�0����7p����F�*>�WB�$1�WUM ��f�s�����y��vs��@
F"�H�`q-I���r���ס����;�2|`[�!5��6���f����0�؈��/�
�~�(�2\���ݤB8�	l��p�����Ϸ|>���y=s�{�YA(S�?���#�J�q�w���|0�#�*�H#O#8�|�������Wx�LH "I�"�~� �PT�GZ�̞P����UU�m�� gϞő#G�#� �v�7����$��BѫV5�nO��\�EH����E|iؔu���J��^�S��uUՐJED��j����ƅ���|��.������oz���<j�f��e(��Fz2u( �B�4d�"d���F�l��62�~�~?��?(u:����s�E��љ�"C
���C@�����$F��<o���jf8C)��HQ��51d��bÉG�d[B���Z7)��m�`��8:�|4���S.B��2+	���i���������^����{�i�g������߾��(d7F�5�W�Ȥ)*�E�T*h6�����@u�)���6@J����.5O�6��6X��$�ܘ��n����C�[>�bP��g-7DKh�S.�J��ȴH��J2��e�(���D�)��F��Κؖ��3��n����TK�>u۲3���$@48�I�`;�i���`�@k	)#0f�iRW�s�kAVgsrr����Y�M\��{��At:����s,F��a²�(��: 4l��Q(I����G�ݍZ��j�&��1��@F}�~����i]υc{x���|gϞM9�����"LLLd�J(<����:����q�E� \
�}����n��iς++����9i�Q��@&���%�U�  8<{�B�.�����,(���􀤮UZ�̃�R��n�C&��F
��jcqq��bjj
ׯ_���\ׅmۉp��Pݧ6ȧp��,..�s��	Sd]YYA��2��V����vq���al�vV$|ݝ{��[,��{�X,��}g�=���#��5"�7o���o���9�����.�p������􏘙9�N$!lqA��`��g��]ם�,�/�&��[��ăY�����F�VC�P2��5K���7g&����O��Ι��JqiwaZ�N�m��{�/�����7>Q9r7}빆gff2����p��MT���6[gt��'�͛�P)�AZ�4����`ȁ8/(d�.����ĤѲ_Y���"fffp��5:tA�b6\�ܐ��2^�A���L;2��.��2��2����+W^�v�~�_�?�)��Ǳ���!�k�Z�z�E4��ϛ��Z�����3���_�"�z����_O�ެ��.���z�*<�G�T�j}*��P+�T*����(ǉ�%]� M,�^7�����ԡ:��������W��u�Ř�M�+�!�ק�i�[W�V��~_�4ߔc�Y�� 3� ��*�E�`K�����w_XX�\�÷��R��F�.?�NdI�Ԓ8����8��&&Է���}0}x�RAp�P�Ԭױ��������_Ǎ7P�T��K/�駟&��Q��W8�nM��(c�E���k�cL3����_>s�|���S�NM���(�J��j}�(�p�ʕ,e}+���ϟ�+���3g� �:-�56J���B� (�v��@������^�U*p-��v�Q�D�1�Pzkyy�ׅB�a'�i�c�4�^*��Rw:Ei����8c�"�����ַ��w�}�/_Nhb�RP��*��+�EQ���j�;p��l[`ee��!�~�<vJJ�0q��	�ˮ�Y������
	0�8תg0�"�J��z��[^�q��q��w�裏"C�>}�|��zrr��֢�n�(���l���ʋ2����Z��N��B4NN(��e#fE1���tb�4�=\%�Ԥ�	%��N�/��ms��LL���7��t�}�����x�wp��a4�M(�2i�����E)^/�Kܬ��/�v'�
�a+ķ��*N�<ER��R
�Xq˲���-8laB�\�|��͛�(��W����u�r�[
@�R}���h��\�\�4���� �5�t��!ͧO�&?��ͽ�����{�M�n�OK;vl���~��������p=a3ġC������{Ϯ{`�R(�h�Z�x�"�~�m\�x1�XB����`�Ǳ�%>���FF�SKI����.\�����-����/��8�>�A�
���S��Ak��@t`��ڇ��W��h�R,CS��L9��*#���h��	萡X,֞x�	r��	���}?��O2ʨ7n�P(d��i+t
�q]7+���a�"����KN���q��1|��� �j�R�T��°�0�cl|���j�ߵq��e���I^ ��b�lC@�`N����'�|���ZCJD��L�;0 P+����?��G�q��*������?�i҇���J�>�u�/}	/��¯_y啇~�����㦅���F��KĂ�z�����_���H�#��{�=��P0Ά>K꒭����׺��H�\9��?\č��8y�q��lG�ȑÀ��	ɼL��� �����[���xZ˄Ӏajj���?���?�����!��j�͘�9fff��\N��_̿g�Px=�{�%�y-�0`T3�\JP��J�B�f��dÄ��g��JШ��\�Q���d�7�����Ɋ�Jg�P��&�/��R�\�Z�dj),	��^�b)�����Xr�9��8�=r�7�n��84ha�L�Px��7��o��/\�����>i��5�ZkQ���y�3����~����g>CZ�V�͒��<Z���Ѥ>qN's�u	�/\Z�9���/cjjՊ/P)�AI�GagV&����%�$}̳ ��G%�V�0p�<QD
��3�Is�!�m۵4)b���ũ�uHڠk�R����z���@޹�w��.°�\׆� F">G�[(��<,wRC���B���&��L���ҥ4��£�^.^�P��O݇˗KX]]I���CBp@3�a4�[7��x���Ą~��73��,�4 �B����
����h�\J�.N�>M]8�5غn!��o��ߧ1����̉� ���;�*��n�!mT��� ������K�"��_�1��r��]�4Ӵ~M �=�K&OAA�E�^P}��p�L�ɥv��Q��Bmo����p=�����m��s�E��scS�%U3�e�l'��m��ia�]��Vy%�m׳q��4>�p
a�s=�}�-��Zkض��}�s��_���͝W4�i
s')P�C值Eݒ�H ��a�0j�.\��R�d���U�Y�~�U���ƛA��j7	X�Q� MR�`� q���6��]�d�+4)(-!���:(
�TJ�����2���	دo7����
�C0�SP������Z��m�s�`=%��p�����{�|��k<˅"b��(�R�D)j*	cX�b���T�� }� �H��+%��.�*Cm�ff�`�_y;BeI�sx�Ǳ��	�������8N�S�?D���>gY ާ  {1D��.k���.@J�w[a׈A���<����"�TԳy˴'F.Ne0�,��7I�)���: h�켛�_��X?������͔a�Bc�2����*�a��צ������9�N[�
tݶ㊬�]ڍ����Ӝ~M�֣)@��DA��p-�vP��K�$��-~��?������`���BufeҮ�j��h�[��(M�.+I��=vy��w~O���JX6�%��7_斯�:$,�!��e.%/���|��S� ,����n@i�ֻ��#�nR�����@(���HH$)F��h��~#�������y$�Cq�� ��i^���v����r6Ob>�W_uC��LG���Y��Јa	aYmȾi�z\8��˧g`�&j q�l�f��dwY�O�����R `d�ڏ��>o;;H#Su�u�h�BMĝ��
C��T�ii�А�}��|��b�Q��~�V��t���	�J�����"�^����7���=/���l���)`u~~�Ւ�k��J�%=�K���,�r^�z�_ovk-L�(H�̸H2Q��1��1�{5�@�5�ޱ�&���O�(Co��o�[��-���]W�ۛ}�����_/������z��]2��h4V��\W �:�g=F�sDG��}dw���3� �Y����d�H�re,;y��=5���hwЈ 8��n��")�\.�ɤ՟�����v��ׂ�"�n�&Hչòh�ä�C���y�T�X\Z�h`k�: 	��6�Kyn�%��<no�,����*��*�h�5H�H����8F pܗG���^�2#�u���{�Y�b��vq������Av�;��\炞m��`�@XQ�5I�˕=��vs�h��Cm439�(���J����&�u=x�kԭ���n�Yc.���zvuu�Q�����N?la%��]�2��ܨ��Hmo�Q�n��h4Ѩ�Q���H�&j����`R{Kd�6l���T��_UkO�0��2� ���]đ��cPm�"��鱁��yTo�G{`<�7£��r	����94��"�� �]�7M�`{!�蹏��j��e���
T(��U?���w�6[_2]V�TL&t�4#�T:���`Ϛ秵�^��v�e��p��w��_��ɣ������.���;�z�Z� 
�F9(�#C�b$�M��n^���c�-D�k�D=f~�"���4{Pđ�6�EQ'�5@�c��&���9f�Tk�m�[�@��d��0Qe�cR=���&���x���\�r)��!�������m�����L�¥��
4i%]������i� ᨔ�ЉL"!�vZ���1˝��^�Q�:m�Rai��F؂�z���z�m��&2����M#�e�����)9ƚ�����0�(�q��: h�Z���l����ʀ�[ǅ 
R�!� �
�T����[�q�ݡdZKPj��#`�H6�'�?�q�:7�>X�ˮ�F�^�x{�I�m�����'e��A�~�C��]]ڣ�I����@k����x�����_k�	Av�6á~rE����T�4��#V��`B����B>�~����\Qj�r�l6�n�q㣏�)�]���5+l�$,��?T��J���g�����N����?�R*x���%8���'O��&8���W��5��͋��N>�弐�3H�j Q����v۝�?��u@
=%R�c��\F�T��xX^ZBP*��h`iyQ'�	���ͲdÕ�f"l��l�h�Z}�h�~��ڰ����),..czz����ZarjZ��햂�z[]��{���[�Ժ	�����ǎ���&�U���Аx�?����G̓�8R��� ���
g� .e��]����C���m4Z-.� �	!A�^���z��f8�6�&�Ţ)Xf���^��5�:0E��կ��
���W05=!,<�У8s�Өպ�����ܰ���X��<0d0�O�b29M	8pl/S������F++�[-�;DF�rv��ZP��h�q��i��s7�Pk4Q�VQ*V�lIt;Aa����7t���/�Ϗ���� �F�g?v��Ҥ�ǐJ����f��(N��90��|��NN�2B��6�s���c���o M�>���~�p�U����`ׄ�#+\J%!8M�bqy	��:��Z��,َ/�����0R+�˘��BE����dO�03zB�\$x���<y�_��>x���cO1��l$q����0q��c��h���U�~	+�&d���%#�7k1*��ɜ%���] ǎ߃��f`���:Ξ=-u	��zd�R�gez�	�hU�n��z/?�w_��&&+F��[�6�&��ܕ��|�)4$���7���p6[ ��?�ۜg��)���x��G0?w�[�]�A�W�9��޺Z �^,���؂\��mw���� RvA�e�\����a��Ӊ���6�V�lЍc8���{��c}��)�u�$NQI	�oY�}�}�-�.�<�.�7�j��H[�)c(ʗ�9�뗯��aձ
J����񅤠@���p�9Un��8n�~��D���*��n�V%.��|�۳8#<0$y���}��^AA�r�<�d���������g��A�삠R��� ���	M�����ӹbñ�?4d�f������|�@���    IEND�B`�PK   sRWZ�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   sRWZ���N/  D&     jsons/user_defined.json�Z�r�F�_�AM�}��Hɖ��mR[*� ��QKFQ���� )�.�Ȯ}���9s��}�����a�'����r������O_����/hB�OV�}t5=���7sw׎��Y3���M�'y]�p�����2�Z7�u3��m��wD'�-V~6-��T�>sJk"�s�(��B޾2^s�}�����UV�f;���o��;��FӜP�Z"d�$�%���;g�
!Y�q\�U�vP���4�$H��^�B ��TAgJ�t7hY�e��'�����X-��Z��LA%�Y���w�����b����c��./�wM] >�z�@�*��]�v�M�
3%x"����buZf��OO�z�[�p�o����=Lg��0/�J$�L����W�l�u�	Z�h�&�|`7��/$ �`���c~>/:𚙄J�ű�rx��J��[j�LX����}>Ƞ��AE }�A2��P�F�� �m(q8@��4?%o.ߒ�A"�!R["�vD���DW�D�Cd�J�0!g���P�!���͈�zD-6$`"I��]io���������&�j�v��<��b>�O]y�x��&ulˠið�G�|{�VG0KzT����O������������������M�+�;����ci����e���X��ί/(�m����]]�T�_�g���{kn�U�.���j��zC��c�]�.k���d|����J��;P�vd8�*}��<� �}�s�/����X��Ň�e��攞����ރO��n19��XM�T����3���5�?�Ge�=ږ�;R�S�d$��Ѧ8H5׌�������UD����%FЌ�����L�'w4��6�&j�#�6H&Z[�
ā'�i��@�DS4S�>h��ws� �(K|�?T�~)��T)#95G��\���S��oO�!�A�W�TG���Q	��k#�%u����j"�OI�%)�s��'�ޣԮ�jr�^M��$i��>'V:JL���G2T�y�8M�V��A
�	�� )��9�62gC�9�dֽ^�Ǫqu���)1������p�ܶ~͗����3&рa\H8����bl&�o��fl&_?4S�T�&��._ʠ��:8n6��ƻ�O�ւW<��[��bw��P��frQ��v�����%zQ0F��2Ԡ��!��s�i��a�V��"��ɻ���>�P�8�ɓ8o�t��9���\qʥ�8u0^`kXO1=J��H}F��[�j
�X,�D�T)�p�N ������&������k�1�z���=���)��%·oT����%�Y|�09fS�1nu`Dd�$i��!3`�*#<^���ۿ���:nO�|]��d~:��pL�f6u�M(z"r!�eR�܃�Un98;4��ƳRmQ$�)�39q�J�[�t�Q�vڸ8p1z���-�7n	W�l� ��v�%{o7-F)����M ��a�&J���=WJ�LZ|�X�9�3T$�S}(�#�B�3�D�9�	���eb��z��?��>P�~�_�?l��M �
|����6�˫��MDoW��눎���W1�\�/c�@�	F�=�\�'���q_�߸6n��GD]�Wp��G���`��oF�����?�<L���&Np�����Ϭ�a?�+hW�&~�pYW�6^LV���0�搓U���Q1Ds'j��SL��O����!&Z�cM䮆!Z����t5�"ˢ��b�����|�'���[����T�x�u��p��=�8�n��m8�����?�a���m�'YA���+��{Ķ_�v5󞌪��0�6�#g�`ǵ0o�PK   sRWZ'.Ǐ�  {�             ��    cirkitFile.jsonPK   sRWZx^��6� _� /           ��  images/00531496-7d3e-47f9-840c-8f79a4e99c6a.pngPK   sRWZWC��)�  � /           ���� images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK   sRWZ��_8
  3
  /           ���{ images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK   sRWZ$���� �� /           ���� images/669aa2f4-fbbf-424d-aa05-a9f27f46a07b.pngPK   sRWZ/�iz$  �$  /           ���i images/750a72b5-fab7-4eeb-bf09-b1fa16e3eb7f.pngPK   sRWZ�Ba�  �  /           ���� images/8da9f3e5-57f2-4cd5-bbab-5c1279684e76.pngPK   sRWZ`$} [ /           ���# images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK   sRWZ� `�5&  0&  /           ��I� images/e181a1ff-876a-43d9-9539-3671c727f4f4.pngPK   sRWZ�E����  :�  /           ���� images/e85fedc0-029f-4b1e-9a1b-73b665cc1a4b.pngPK   sRWZ�+�s;  z;  /           ���g images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK   sRWZ���N/  D&             ��j� jsons/user_defined.jsonPK      $  Ϊ   